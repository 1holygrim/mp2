XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�� �ggr{)������ި}ֿ���.5j�\�x�>���<��� _҆ZL���\={t�)@�Or�9s z�� ���RKo�ڬ� U�yc���]*<�i!vݞܟ &����DعjNU�Sk�'�U�9Bt|����k g������ku�魼P{��g�@&X�����E�j^�(��E���!�T���ޛ�$G~���4���
�;Ȳ����;?]]2����ܼ/f�OjtK�Sts$O;]9h���]��-���.P��E�ן�T0	���ƥ�U˿F=ˠ�0ńѢ�X��m��7�i�U!��c�#^�,��= A/'P�#͉�}��64c����)S��4�'.���I�k�L�#�J���w+�ϳ��]3&�b
�7lt�keCn'�βY��(<*�o�B���g���GK��T#g� ���1��b�T9Y&��@�q�r�ݼI$�M?10�j�E��A�����?�Z`�..�b�DL����*)㜬8Ҍ'�܉�J��)����!~~ףo���n���!2{���0��Co�+`�S�2F���ek�Ǆ�̵�eZO�o"ˏj)���DL�:�md��O����'�ǱM٬|pT��K�[�ǚB��s
r.JL�!_���n&����S�0��"F+��\���酮�7X���,���(�C��R/n�
"��]x�o��0F,�>� ��R�{Q�-Dd��c��c��qazP{4�C��f��8�XlxVHYEB    dd8f    2160V��������J����lګS��+|nJ)��#��j	��mߧ܁"����8��>�t��ގ�6�c�u�ͺ쌍?�FD#�;�u���Q��|+J�E�K��LNi�Ar0�U�i�s^/�ۺ�ߏ��o�P�.HF�_Z��E�a��Y��,'�j:p��<ʹB� �vZKQ
!E{��nE40��Ӹ���杼��u�Y=]��!V~�ý��2�w�����F��t2it�zP�yr�?IzX@F��T�tla��l�\�ᾄO���C��e=�uIsz�N��y�/IC-1ZH��}���Ŀ�)?�V��~�f�d@y��
�����*l}}�r{�H��_�b�b�C� o'��˶��$H�oUy$�u�ݤ<����ov���&l�a���C+Dd_��N�1�ʖ5��r�W��]冖�0P���jc�`Ab�Iz�ۜ�x�j��γ��}�
����a��ڍ�2}���w���t>u���r5�pl�"��Z���(c�WoX6�1.�k�� ��"�m�_�d�h�H�-��9�p�g�T���K������2�捪^g�3�CC`<S� 2�����7(���&Ƞ]J���WҙJ ���=Pc���|F)}L]�4уOi�L���ћ|DVay�G6o������[��vN�P`dR�/wƱ�� ���>��̖Y���ms���ӫ��IL[l���0rfi��) �m/��V("BVGmu�� ^���%����;��T��G��A������a��YE��4��GS�V��u����I1��b��$�[��d���ͨ+�KK�{o��\P-��a�c���4d��E�̠@�kz;e�*���M���[��i�fTK�VLx�B�qkk�����ig{�Xk9�3�'X�3�V������4��dUt�^��_�..ki�c��5�G=H^����r^���+1a��6�ҀyăÃ��Y�q$�>�g���=x�'����}�s�)�6a�:�:����e����+et�G1����������_|���=�1r1A(��(���MG@6���I9G��&��7�g��{�;���»?gF����Po~�i�2Ţ9(G���6�߁�H������>Ss;ee?�+�CS�s��T�]�O�?s�S��k��׊J+B��*G�"���� f/��t�N��H�r��fB�K�;U�d>Hf�t^�h���v��B�Π�E{m�`^������Ɯ�x��|����Ye	b�  �-������&����w�O�ڃ����/^1�%0Q���w�(m��/�˸-~������9�{�ֶ�T����M,���.c2�B���U9G�߷�OZ�2m��y����]��O�:����Ι�И�]�f`�����C����K�{�����c�>�x�L\��RU�u��r8�d�b��ۓ>�c�F��W�2���1�'BG�a�����6Do���U.��d���+q(NQO��慇7�Sw������h���AT�@��hӚ-q.6}����@��s��û����������w��(6�$��x3�J	�}?.�hS���"	b�8��b���A�r��Ь��w�lqx����\(2+�R���s4{{&*1uΚ��Á;])�O��u:A�X��ư��g�`i�n�H2��,�y�S���A��7�k\#)c�b����dPF��� *��;����F��&��"��pܤQ&��u�)���;_ï�w}�>�)��1G;<Cބ^ބ�~�?޼	�#�߽�Dü�ҥ���=r�����}��n�b�(d�		KϽk_��>J�+\��N� "�Y\��>r�eG�~��M[���.�ƻ׬�qj��la�dJg%f؄u����箻h�B�h11uǖ���j�5�$�p�k��C��`uZ��{����6x�����%@&�
���+�z|11�Ke@ �g��T�X����������V$&]K�D� ���
;��2��yt@ك�	4��۝������ϓ��'�XF��
J	���oY�Zv�+'t5�!�2�ΫpDY&^kn��Y�FX|w�|0|�{4Gu-�@�.���4�U;�ϕ�*e�c��g���?y=�ݒ�����(΄X�{� �bzr��16����,�l�v�<�6��j �;"��y����k��wG��j�6�m~��69OhNU�-�
g�|�&���t*�d��j��N&� ��S���%uuDU������@������xŅ���7�+��rBP67���{���/!��V_��i���00������=Z�]�g�L�$wT��K����C��l����W������AEyjwZ��Ps\���c�(�T��_$�Ԧ�m��R\�����8� �'O�uivկ���(V~�+hر]���ǴOFYg("%OVG0Ӱp8ܗ�k@�;���G@���d�:��<�eoq�V�4�XǊ�fz���\����E;���oY2@hUDS�D�<�[�|0k��B=K�!EY�ش��cv0_�0�A���ղ'U���˚�
� @j
�Y��#?#m7cVbG���Z�g9��3����߾Y$OQ#p�C1D�D�R��oku�o��^�ɂ�R�N�°�9����~��/lmwS�t��r"ǻҞh��+mV���P�{���<�+�6���Zw�[�w�5Y*��%(�IЦEW�C��쉡��9���1��g�����B� U�FlWn�s���K��C}3/9���m�}�q~=TC�D����Mh$����pn�ys$��b�d���>?�_@{5Ԍt��x0����`�rW�w����wH���pya@���Ä �X����o�\M�=��k������}�{�XPc{��zR6j�b�ל�)
l�j儲t�Q�y��V��=��v���Y�\����@<��At\�f�1x�[1 6��SY1�M1�6FL���Ь��KB���1p|D�ƚ"�df/�I��0 ES^�-D:T�<{J��\��Q��/����y�Q(6f�p�8�H�<�[-�^�6���b��]����M�JfL��{�iha�A�_$B��G'��};5�_D�	�BDd��j�[r�d�J�X�0�y@d��_[�w3���*xz�OP=��}3O,�ٚw�����*U����/\O��:.��|���yݶI4��7�T���X�X3A������
E�l��N����գ�7I6��&�fB��W�������ք�g.))��ב|j4B����iwq��jH����A}S���A4Ox��1�u,vںӣ�&n�JR]L�1�ꧭ ��$2����]j���ʻ���͍aU;.<љ�N�ߗ(!-�jA��L&!,.�>Dw���]�b�p�A2%�ɺ}A�o�5W3#6?k0TẀ��Ȳp��c掊��mw���Ҕ�^\Fw�2�B��<Ϋ'ms�Op?��T{��fUֻ�Y⩐d� P%�,DR�\R��6-	Ɖ��I�UO�9�w�y�, ��!�ʈʦ�#`��x�=ʆ\��7��P4�>������GLR�s��Hy)!*I��Y�AR#�s��$�Osیʞ&��L(Қ
�"�:x���B�1E���M/B�$�f%t��K�Zrz�[�i|O0韕�('���ޫ6<4.ҹ����0���T������L����n�~�N�I��u\f嵙W�����0���(O�1��bQ��Jj�܋�b���ů�ܭ7F�;	�[pܱz另��r�J�p�����襭%�ܴ����'�N�E:L�Z�դ�%�e������vR+ߗ}����wp�iד�%s�Wo6K���h��3X���S��i�C�����^-�xK�f�i�eI~��zu���IJ�53S��y����FK:�w�&�k����n2��O��GJ�C]y�1��SU$���]F����U�#Q7�1n����g� �
�.��Ĩ����	�������F:=Q� ���|'��Fq-�m�SQ �Ns�3>�����#�&������ׯzs��w���s� ����Q`����~�<��3�v�F�Y�q��5���=�B��F�?d����O4.�O�sO�Pw�>�����rZ��d��^�!ˎe�4=-n�to�!EJl�$n���k�u�TL�1���v��siY<|Վw�5�4HA���u}�7lV��j�%�y��|{��Fa¦)M'lWQ�o4� vw�A��7٥܉Dr�
����}x��m��H�X�� ���Ig���m�9G�dl�" B��[z��7&�����{)oa,��]��-,�w�H4x�D2}��i���� Vm�y��
~��a�A�N�!��������q�^�e*~p
l�t� ������VM��ib���;͞'Q,��΂��<�I�@z�a*��V�$ka�F9��3�5JM[���s�,�A,��[�A��8Ӗ����k�������A%"�ޟ�)����!Z�9y��D��������e�H��ᱞobO�7nVW�� &wB�܍�����HD���@G��k����X�5�`��b�|�և��C�Fc����z+a^՛�Y���u6˸�R�pm��Y���a��!��|��JT�T1�փ������R����%��� �|0��ǯ8��=���:����;���$m���E�����wel|Ԃ�<��Er��B�p�u��0�"�AC��1�Z$� �{�X�:���z�.��gifSnP9^�#@	l?[�Y`��Ty�~iz'���M�ɑEP
�*���r�{J���c��g�s��e�7�8c�'n��o�Ǭ6P}�W��v�K�"+�)~e�Y`Ln)�]g��4R�:��z�-�.�lj�4�s��.�*m�ñE��۠�����{2K?^�%ģ��v٦�j����W����A��W9§�* LwJ����0%�$|S�L��1Ȃ*~�����ȟz���%�~b��y��1i��w�9kj�Q�'��e7���s��BH���I9L �?PJ�ӱ�@,ds��� ����88˄��]5��5�R*��$��I����ݼ����܋���fN��`C��[�d�`�z��F�S����M�i�
G����tV�x� 	�E��;� �qA~^`��Y���x�e��#�*F�yc��)c�����b���B�,,
_�B�1��� �hE�u�5\�@p��Q�m��*�f3Tr�����՗��EkR�.nX\1)��m���^̻%�k1N��X$�7T���g�ް�aO<1g��OC����·�q6T6Y�6��^�aז�%S�gZ�;I��7 ���d�@�Y����YT�!��������T�F9ƻ��^��`
�����!�r�[�&t / ����o@���J}y+U>�MձFڵCW1)iT�װ��(����`.y9�'�nw�P��
��ô�O?��0y9�'|��(�:,:e�S)T��+��g���.�Iߥ���֖�?h��"���{�-�qwA��j��oU��z�G��A5�\�3�����	�z��~%m��	<���?�S�3��-��ZվHq�o�G�����&1���9��2	ҷ׬`i_ꄻ|�d�Z��Urû�P�3dZ1�����b^��+O<���4��b�x�!l���P {��i�6~�k�6�_��d�z��!'uj�+!�0��� eR��T4�U����DNo��N�(�I�D�b�Q��V}�xx���ԙ��[�����;��O'f�6�)�򫎲A��y��+�&޸�9O�s�B6��m'%
�,k��>��;Su���
�v��UK�cb4��(pS��w(�@SqǏ>N��#�[m�?,��ǜF�K;�5��>�{R$��TNn:����]��qu�Jl���B�N� 0�M�e���P|����]�
Cz:�$I
�s�9���>�f�ϛa�ܩ8�BD���ţ����h����B�;3HJK�z��I�J�',�1K����x��� +���륶�E����|����
��~�ԦV�X���ca�C���PGr�h~�C��%$xC�˙!a�_q��������(��R]�t�ܜ{0�~�O�3���!7UW'��Þ�}�S��RQ��D=��Ճ��ͫ��ϒ�{��)YCUN��3t�~��D�镬^�%v�-�Q�}�5.,̳'6X���;�Q�����Vi���\�8���-C_�P�Z�������f�T��4��/��r�S���@��p�2�̛��^�k�9K���cx��E�ڰ?�������zz�e?������͚O���d�bK���U��3���PF�]��5��2����{�ȍ2�
-�eڒ��7���vaD���cV�Վ�W��ƽ&ڜv��Fg���)�r���s��P��oVä￼{Db�4!sd��<
+[AP��f>a�6���~M'\g��)�h{e�|�M+j8+.�&Z����:�,��	�)�"d)X!��.w&±еiSw{02i~Z̘8a�qOmǥ[��Bf�N�gd�"�l"�.�G�E*�#�ȣ*`�ӧ���k�����6_bY�[kbi���_��wj��?�79�?�DD\�t�c�ys@�ܲ�|���O�e}�Iu�y��������,�ʢbp�6�'�9R�rps����-���%�m�]h�qZ�ق�dv�_Hb�k/8���~ݹ��o�KF�����U�;��qXq�;f����2���3��x&T��:��Y������`�M��{��1��C�\N'P2�Q �(��+l���5Ŕ1Z�G���kL�4Q-J�6ҷ�u	�sB�B;�*U�:o�b�Cِ�c����ժ&7�"e<�`;��	eGUDEr��|����a�~2x�_N� ��[�q��y��8�r����י��z5�����68D�����$�&0�)��7.��d�q{Qt�@�����j����
Q��I�&=����:׸d�	��{gq}0qpc�����d���#I�a�������p	��ݚ��m
�-�?�؇.<��M�F�3"��*��hp.`�Dl�¤�7}3lx��|��7�� �&#�
&�I֩٣�w��H��i(_oo�~�`�1I���+R��Dj��1����L꟫Y� :z+r³=����.��*��2�cH2����l��sc+/c�P��G���:���YG��Cq�	%@zh�D����H�D"ˡ�)4�t����Q���O,tڏF�v,��B�8*
�F�n�����۠��77��?�sc��9϶_�[ǽ�(R�۠~{�Uʫ��� �Ŭ�3Ì����q��y&�M@���YT�fl�U9@����܍t&79C��`7}vh�0��h���iI���:�aڢj��=�ޒL�'��x�IGnD��M�aS�Kz�&��5�3)a�����:�ׇM�DψJ&y�7����co�\m3{f��a ��ކ~@fg'bD�@{u���P�/e�끩�n`m���[�׎.s~aO&��C"7�s�	�'iQFbD-�
�F[V��&��jZ�����c���s)#�
,l[M�[�����c�Eｐ:R��O�̛��bx��ٟ�2�G����b�w�62���f�(
������4չs����������h�[��-[]9�"��?�K��{n���p�h<^���D~>#����o���`����֨/�H��Z;b���&M�+��%��6S�4-_(#f���z\�iA	C��&Ary�.�g�|(�6/�ä ��w٧t�	ǖ�����t�t@&��ss�����F�t�d6e:xkZT	�~�����F�uJ1�3�nϏ=$�Snx�����PU�^P	���׍_��JG��>c��]��՚�2��MH-��c�_�C(�z^T/;ե1�H;���)�úٯc��M��8��vBO~�N�љQ���|�K������Z3��į�ӫKY����;r*5w�6~]$��_��p+��d�>���fo�|����[~&(D&�m�t�ߋ ���Z_�9�Y����{������_�ۍ�-��@����
��lۊow���r[�0�6������4���`�>�IQU�	���̢��}Ǿt�_V$���[�JI3��x�w��&���s;������]v�űmzǢ+�j�BC��3$�u�æ�9�r)H^��tb�T�Ŝ-�h��D�m*6��("�f�ܯ��.�߰�b]���<7�_���2�O0Lm:W�W��i��=z<�������<
�2�{�x�q�/�Ҍbjջ
͚|�~w>w�n|0g�=o�ź�َ�n� �	���3�_�gH�p'ﶠ�w�{Mx���