XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��T�ZO��x 6�w�������A蜻���"��
�S�+ʚ~2G-�f_�E�2&�{��9 ���_�>y���d�P����YI�4���MK��l�m~�N;�t%�}�"x�&���d,q�3���#X[�)�8B\�� ����j���������1h�K�	�	+�C� ��ȽົxLM>ÚЧE{� ��Ld�>��Vh�8n�k'�P�DV~UH<���%��s�C�����5��)���DD�&I �s,������Ŷ#c��Rq�1�n�H�[݂y���P�2�@S�Hs���O�#xj�'R�(��*�qQ]A��*��P�WM�rN�PԾ:	���cxq+c[IK�Fy$&|�q��Ĭ웞F/jc�`�"MH~3�;�Z-u��Wd�Ћze�����s�H�E���-!�3x��:�*SvJJYrH����h�VeXZ�~R��Aw��̅�_��n��Z'������2��./�&��!=Y ����fs����ܬ78)rZ.�C��������������w�@� ���(�(�-]~�먬�^���s�L&��;9�<F�uUz�i��G��B���B��͈^�ʨs`���{Ym��(�Ѣ�Ka���"�K�K����ˉ��Z�h������jK�xRM�����WUIWQ@M憺���ϬY�c��ϲ�{�eL=�Z��w���h��S�m��w{2F��?��#���en6�0�d�c��"��L�w�Ho�O�	�?�yJ�G Mc�Ng:ʹ��he��l�XlxVHYEB    1853     810������{�qH�A����g^l� �B��T(��S�H@4���g!��$�E�b�6{3r8����W�P(޽<P���y��7gq����Be"� h.H�o}3;8���׫�Do��I�AE��"�l� �#<WN�C��`Ksi��]��� P�KG�Y��/�t�H~�e�D���T���S�����5^īR\0���D����|��Xu���F4�-��T�a���TG�UhS=�B7��'Zs�:�ݐ�T�e��5�UɐD�j[�?�Ѹ����m��E"qlA�2IT]s٭1Z�\f�N��Z�=Wd�]�I�����}��u����nKS�} L$oԚ��������B"�5�lZMf��*����<DR
�2_��XE�D��zZ�hI	A�� ���#9�>#�l������o񲙻2@�5(��.���kdn���*xU8$�p�ڥ����N���o�y3���.h�wƂ"Y�����3���g~N��6=�I�X�3�����I��ҫ�J���>/�Qh���<j�
q���yN��	m��X�#��W#�}&vj�ؒػ�`O�]6���B�'�o}�c��9�!|9`���1�[PwQ��M��JHL���siՂ��~S�G&_��7CUXx���(6��(hyK��!��g�o��-��x��N_��sy���Fg����r7�I���{�W���2e�5n�7��%�f����8��Plܿ����!�Lf3̐m�_�͔�����[؜�3���s\��}]�8����������/��0���3��5�5���,y#���;U��}]�5j3�y�M�ӓ2�7��\UoM��Q��7m�E�ڝ #>� �m��D�����ED���r�����������6����cf�#��9�h�v��v���-�(�c�%��ݢ��я)���V��Ş�C�5y���F������Dv���PY��a������qTO��_.	�����Ԓ5��%9�wtp�,�כ�_�y����0�H���s�H���ߠ����|B��l�:���s�o�{E�u�Ÿ!���UF�8&���Iq�����a��Z�sS���E[t��xʒ��/-�IT� ��×>fqZ��]jP��w��_9M�C�q�N�����Ө�<D�6)���/�}�o +RpQt�L27 4\��Dj�^랡}��u�)K�m��Ⱥ�D�WY��qE��'i�3�
�*����X�|c"�,�Ii8|K���	n�#s-��v���y$�Cug��Ƴ�o����.�'Q	.!��+E��1�tS��+9_L�'�YW$�J3  � � �&���x��+)%�(�}]�?�3in�wz(~�+�@�\ఢUkFݒ))b�A�juy�5q������y�HdA-�z���y�.!'�e���n˯�o�q]fF>�������I7�y��ղ\M$·�g�tB	'i_�K��n�oY��%���g�kyp_is�G���2JxER���T�5n����=�p���.��<�wjX-f4 12O߬�Ӣn�8<�v�*N>��a���anw;��孱@���q��d#Ԅ̯�DB	abPi}NGw�h�:�#����3�-7֙�g�4�W㵙�������άyu�z(F��`��O��J�+'�Q��s�,�n�����tՙ�j?i���p`����@N�][ڬM�,�a7����K�Er��ٞU�c��u���ئl.vs;���uG�����|�Qr��R��6��8 \��n+/�6����õ�[��'���H'���"�O�0=/Ƅn�SU�]!����k��qqp�kLK�\uZ!��'W�0a�:�#yDVAe�X��}�#5��W/�8$�q��gY����� &��wAJC��Y&nXn/�t���s��AǑX����:TO��n���A�^p�G2;��%�X[�C�#���T�G�����%����:(��D��!	�M:�n<������ug9%I���l��K�O2"�ԛ%�qx��tS�