XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��.��bD�R�D��XY`���K���J�������>�K�����;���z���8S(�j�Y;���
J�e�*�;��
^�A��Q��1��C�Ç���1��t���S%���i*�g\��}��'��7@u��Eж��?�.3��:-�@c�BOf��� ����br�=��#��ͦU�X56�g�a}�����.8�F���<�j�6�8�v)Q��A:�ʇ�7�~����phUN��,�+~]�<�Z$�����oπW,�ɛg�{K����;,A975[&��CV{�������nB,�zg�q���G���|��$�'��蠙�E�3� ��	6��I����1C ��haP|�������fO>譓�Y9OI�����m�
��E��[����Ck9��%�-氯�T�;FD*#ƿ��+ˣ��Q�t����ː�î,:a��~��~���ԭ��Љ;� ��Qt$�5���6�M~��>�fRZp��y,J`�E@{��k�AK��ee�zkL2��F����v%$���&�7_��Pf�煐G!2��VG�Ԕd��^�-�m�Zk ��50[5���h����9�~: rh��IQ��l���� ���:��]w�LT�1{��=���')K�X���Z����$˻-������ ����ry��л��4묀�Q5�&ŉ>��lyR���������Z�!yղpCT3D�Z���(�)�I��Ǝ��Jյ`w��YѩuOI���LV�L�h��!�XlxVHYEB    fa00    1f10�!����ɟ��hX�ja�Y�LMMƃ�dw�Z�F���rO4(5���qxM�J��`�.@��*Օދ~dc�����=�F�۾Gn�8�R>,�@�)��)��c�W�|����$s\z����*q���3&n������M2ת�A��g��<TgEVZ��p�0j��� �oW��Ev�8�e�a��*�M	{��g��h�}��$�zɉsb(��ã�o���  ��!G��+����a~�$��#=�n���z�#g
�zC��N/���X8o�{87�Gus9��/���L�f��+
�t�5��sm�9������j+ZN_��u�PO���bQ=sJPא��fX|l��L`�?���2�tNv@��ۚ�R'�&�8��6a����lJ���[-X�,�9���N�k���Bp;f.���3�Q�$���DS��/���=+:M��0�~��l�w�����P��a/*�D6�W�8�T�XRl"��z��kս��K�B��}��3l�r�����@��Oq�TK��楫)_�ޜ�֕���`l�8���	`���xxR�i������9 �۫�c^U*���t�1��d^���<oW�YK�%>om,*�z����<��L�x���a�a/=�]X����a� �U2��|8
�V	;�T?!��;��;sm17fv� c�9�z�US³ѧ���Zs���w�8���KВx�;�J��in���G���#�gj.m���:�<FQߩ��*�h"d�|�G��F������k�*����+���T'�E��NQʧsJ�8ծm�o��=Ă��#�iF7�2$tX��;&�UOF.U�w/j��GD�2����	l�,g�_R�6��3oW����Zb	��ɫ�EE|3�E��JY���X4E���P��$�P��>1X���l��\�K2��^�Gr{0b"��}{���r�7�>��Ơ�����CR������ /O���]�]��Oyr��c���65%��_�IRB�/�N��-I�uFS'�����>�]�)x�qS��S͎>�6B�kT58C4]�YM'��t8;��i��.�
h?�/�ǁ5�8}yR���w���.s]�:H0����Pq���'�L��e�ͩ�6gBpe���cɋ��4;�'��m�}>�|��"d�"�R;�l��[�8*��b�F��513ҙ@���ۥ�n��O~��{�^@:C}.��ekښ{x��H3E:��^�3аg�ƀe
SΜL�9j�\x'�ES�?&{���� _��mVoC�9E�]����@��(ץ�E0�
�G�.ڝ&7~���	.>�B��R*u�fNz�@}�˔�4�q�|�|f7��H��0@�b�I��P븧��+E6���@�e�û(z��:�x�!�������{C����R�c��FC��	��eR!$ �H*�Y�3a��H[)A��B�X��Utb�I���Cg�?JY�:^�Qr0t�#��9�}�t�!�]�k��Q�GuN���)���$\�q�7�[�{�J�����ʑ�cd�'`g:��В���4�mI��)D�9��U�ޣ�G]�m�<�X� �b�9��c'o�q)���,�VD����/H�mkxkLq�&��AQ��w�l=r��A^B�W�)�W���i�5��VR��������U��cB�b��@Xdk�4�w4��]��%�u�L�uq}��5��W��d%�)��fK�Am�?���gl�h<��*�������ك�l[����d�g
,g��Ƭq,Jڒ���<�V��AO�0M* jݎv�*�0���>�v�GT�%�� �F�f#:׏
l�4'�����Ec ��]�ih�1�{>�����1����#Fih�c=e��_�j�dG׹��{Y^�N��I�\���nk�O�D$�Bt=|�:����O��`�d����xJ��, ����J�患�*��p#��Q�,"^��qj�t,��k.�I����Q����m��+�E���Q��}�Y\�}�m��k��J߸�W`�d5v:����Y鶇H�&���ID�X�e��A�}���Ŗbv��BS�D��D�-���.��/I9yLDQ�'��d��@�&F�DE"/�G�6O���;w70-3��m%1;;Q�zF*iɆtFT�c�"�yY�l��|
��m�����b���4��r�5rA(/��2�Ԥ���|w+uj􂟐���؅m��e���\�c���r��ga�^*T��N���QT</���=���|6�!'4mc��.��́=6�� �u�W1ֺRkQS���0���h� s����9.���<�vvp�P��8��m �ZJb8Pm*�j캇"Xr�c5�����P�G�0	�g�1�زZJ�����-q6�It�ю�(�x��cc�������ȧ�ٓb7�BRZ���Z��x�z�b����@�UP	�,�2����0[���Z��l�1�޲����t���J/��S�4H }]B��|~�B�D�C3K%$)l&�*Y�w,9���8|��7�`���'�=+Fp��V���w9^�g+L�7M�YM+�l��eB�;^K�V0uu�M��F�+��@�xD�i�24�i)�i)G���*ki�c�mz��K�A~�ۖ��[J7yz�a���+�d:�q�bA����h�u����<3u����91�Y'K%����Ho�:q%@+��I#�x/B��O�J�y?�\yfߵ#r�Z6: �R������S�UR�4��	]��^	�X�P�S�$�{�P�
X�r����|��q溻���'s�����P���q�`�	��N��O3a�~����*�Agna$�z�|�Z�\4U���E ���0l�M	�\}d�7Ao��%�0���|��g��C\��6]b^��~��إi<����>oq��4Ѱ��Ѓ�}=j=9�Ze��TC�pNAnĔ~ir^J���(#�����)s�S�����¨����fn����GTa�?���t�Z`\xUsT���X�%5��b��%��ʙ��~�۠Z�>��T���2fFB^|>J��z��� ����@�)Q�I����ۄ�\������ܵ���,�0��0����?;sm�-A��@�1�"�$8@�9yL���%���?L;�ǩ���*,i����벒�Ǉ;�K�dá�Fk�*�RL.%�Kj��qi�U�O�a
�/l������@�rO�v�/�O(D��CaK�[���M��Y�M�P���SU)տ�e�>�����}���άC��R[y#�I�wŤ���_A��G��T��s\�P��s�q��ܹ�E�"��PDM���y��t�Ӳ0)P�OL"�ҿo�ZN�f�f����䂻�O�叔ZI�G��r�S	��H�����j�j��@�3�8 ���xLay�v���ㇴֹĜ�)L�a/Ց���n���(�u�OI��1�6�4��ta0��o0�jO���1��e�ᙄ8��e?�O�'H�y��+Q0��Ԋ���`p�b���m��;<c8#T��+_��W-6ww@�5���q��m�.�
vЇ$�E	Hy�β�RYކ�˧ ��kָ�s\7�p��w��6�����%�Bs��^V�,X
��z���=�-��$�~��Y������s�!�q ��P��n�\Ǉ���-Fk�̞uӍ��O̊i倨a[����=��;��k��p?~]�%�#y���xM5��o��r?��t���ge�����S�tw�������,�>�o6#��������:SG��23.���ӥn;��0:�6�2��A���T�
����a�dҲ#m��ذﶕK8H�9�q��J/i�h'��� �� �VQ'.���P��0fJ�A�nn�c>H��x������s��GN�T3�j6ǡ���1ǃ���zEJ6ي*;\/=�9mk��4�É�r����Nwp�(By@>Ps/ӡ�����o��	$�����OU~(����Bc��c�?���RM���/�K�9���"�й[����̇Gc6E�-K٤ʃ}
?7%J:����h����A���0�S�#�~U�9Ҵb�c�A~��_�����,�9�������by	Հ]����;���O�4��)���Pň2�"���8t�ʟ��nM�5ئ�R%B�i�V�淍�L1�>���W�AWM�.dn�$g�v���G���"��í�yp�]�ږ�U�c������<r�Se�u-և���$��\p9�<�V*��V���ِ/�Y�JJ��M~�s���)�Ҫ��$�������V�����w�&���Me=#ٗ��$�
r?�vh@��jbM��|ڇU<{�$F����$����FR'���]<S���ڄa\����i�8aF�l�N�jպ�禛�g��Vヾ�
�dR3�rw����t$&'m��vX޳���I!p��ˏ��Qc�ڙ+:�E��������d7� �e���8%V��B�S��e!���?S�\����c"��5����߭k��谴��PpT*U�g�Dۈ��iF��$�����|.�V���e���p�n4����n-�mwx�[~���=S�:V��Pj��w�z<dk�\O�8T��ks�V��(���m��D\C
*Gk�x�dc���שSn�@���K�wz�Q�1=�2��k�9t�;�E;h-�_���^(�|�νX����ax����*�XF�]rPQdz?�ff�V�8�0�Z���i@�ɞ)��!/���%��E�I�h+�9�T��m<*m��g�R��eCg_R3)�3��F��-�u1iC��lšROq	=8#v"��v�����z������K[�3����
�ŧ�ď@�ʣ��=$ �*����Da�|i"Wla�����^�-�O��!���шyD�>J����[BU���I�=�,7	�{
j2�4�q�j��J 9 �~G�	��-�ǐP�cG'��
^YKVʛ}���q�@��9Գ#�q�E��*�����>�S���Jq�~1���%r���m���E2�!�1��]&�\�(a��JJJ�:N���yJ� eL�|/`gx�}�g,�`������m	��8�/i��L���*�|�e�P��l�f8c,J�BN����J�/���=��s��u��2� I�E��y��E�Ao��-{Y�`��y�YK��r�~�U�!��� �cR�$^�G��sC����Ф��fd5��o���P��ىQ۬�I���c2���M�f+�YΤ����+.[8���]��l5�1n���e���cW��(��-r�
�����̳�D���<�l��������ͳ�eg_�����_���|༹�0$F�@��k��t�e�����&�t��<���G�S<��V���<�>��(�6	f��Q���U����/r��j�یT*D˱^�VB�i!J��`,S���߹l}�ź�=�=�����"Q�Rb�F$_��	�wRb6�����ˣ�������vKv���f�+�V�Â%���c��Zc����L7�i�{&�5�^N��6��$c�_w��`���9'�5X�#>�U�W'6�N8����ڀʪ�~*_E+G�;j/ΓR��=)XK�/�nW��e�'��;�#�21N�Jo����$V���a3������#׈�TM��jN��h[�@v	���x��Ca����a�����o=$'*�:�H�Q��޲LS�R������;'g�Ǐ���hE~�޲,�
ݯ(}�l9ʄtg�(�n����?(ji�����&����F�5��-�V2W
�ƅb5�36��M�X�]t����cZ4�}H��7�Ԥ�m���R0��j�_��t�ᄜu�
;��c4n7O\@
�P�-��{25�x�$]=z��������P�:���'@�b3�	t��2��Ĭ�L����,�4����ͬC�/�u$�P]��zk���/l��� �����t��4 �ܲ���y�Ch�tV#����I}�NyZ�< ���Ń0�L&�����2���Jh���@�1%�$���Ʈ�O�A�#/	C��*�|n��g����zi!w�L�	2��T�vؘU��Շ�V���J��$R�5dRFj��Wj���v]?os%�P(}��I�Ie����J8�v��z���s]4� ��C�J`�"ɑR+�%�kȑ��N�Pg��V$�(ݎ;+K��X1	�/['��Tڱ���6�C��vf�# �H��Z��mR �d��gZqx�\�?jMe��ߣ�)�֐O$��]�%�����rKV����cdH$qO�e�nB��������G��[�z)y��ۍ���w|��"�<&�[��m�}�d�B�d_l�3�]��J`�J�3D���4��QbE!u�y�`�WX�I�*��ؓ��]cN�@�I�%G�玁�����&�SV��� xl\���ݳX>�Q��#	�K#i�5�3�F�>��+�2�����K#0o���7Ȍ�M���}U�B��o���%�*����k����U�5��`����Zk�ؘ�(x�V���z��O�Y����%:
jn8���ǵi��_α�����1����۽�ۅ8�����A[q��5�4��g�Aic��p"�����rq*<�Kk~�5j�B�Ȱ������p���N��#�7��Ơ;����y��1��
]�W��7�:��<�+ �	��?�kK$ P	X����Q�0U�i�]��O��YՔ��X�;����'�.r��ډ8 tܭ�!VZm�6݄r���ɼ�c�����)�r:f<�c;�d��\�!3���X�^��)�!|�W�Ě坈}(�),>���:%��+���[����Gr\��`��q�95P���	�6?��_�E�?|��eY���Oo<��Jc��#(T�$�e�20�E����6m�˰~��J�qYr�qi��Y-~����������IP�VK��uN�%�:k�u.#�ν;��x��R��� ٺ(�j�>�N����^�N����}K��F�x�ݬ��&��Ȱ�����=�I���h&�Wն�4�$�x�����f@Z����T�����m�!-��Ć3�5�A=x;��%Z���J�������!-v��}�a��� �R��ї��9Q�Y�_�bҭ�#�e�w&Rq(Lv�K�8�Ox��# ��ѹ��H��ڶ}�y}ӬT��:P���[��x����"i��40㰫������}w�#Fe#�yB!�b�r�+ҵ
9(o��J�9І�<��$�X��, �hQ���.!��\Ĥ
8s�h�7��Ӻ˫F`s�w����dv�>{�A8�Z3ox�WP�~�TO8������X����̝��֡�5�+���[���l�?�(,'�߷=���Y��y)o`r���
ޘ��W�t?�X�\�%�zd��֦�'}���%#�_@��'6�C�W����=��+��$jD�m�����zg���T @�]�2; D���L��?�\����pg��Qs���e2���q���݉_37�����K��l������HH��A���]��~���]�t��~P�`�'��E��lb~�_��9'x�h�G����É��;Z�L�^ӢL,����6ً���%��_cAU��a�l���ҋ����ac��>�/�ъM�Ҥ�|�� ������f7 �*�_����ƄW�u���JNW�v*oE�x'g
�j�p� �51^ݽ��R���c����s�M���\$�@�f؛n�T�HΑ�+s�B�&��I���o#u���2�
Zq��
)XqXlxVHYEB    db34    23b0Ҝ\� R��7�d���u
NQ�y�Ƀ���oEP0�&��t�oK�&�,�F�QQ�NO�S�QB	bҒ��Z%a�xw�Z��33xNT%��(��N��j�?�Ƶ�i�Yc�-�D�!�����YC�z�3��>���xO�tk��Wlg���9=�A���ťhKa7�V�5E1 �9�W6�X ��d/R�nS���������f��͎�M�{�e�mx��xܾ����%Man�yl���8m����������\�Q�@��)�Z2��T�b�u� ktQ��0^�0�I�k �p��E�r%[YR�tc� ���}"\�gy=b2�MS%;��!a ��z�H�I��.���O��3�����[
ԭ���1�ۻ���t�Q�x�4� H�(��*�U�<Ɏы�]h�k>���r);Qo��x�Ѡ����X��l���T;�%T��흫`YR���/��#�0�Hyʦ�~��%I]�/3�P0��g$_}!���.٭}�p`�����@�5O�v�e�m�`Ip_���0�^XR�g$�y��@K��Y%.�}�kt�>�P��鯠�jum��0	E�s��٧�GR����1�����rF�v�)n�7�ζ�3qD�畖n:�:�t�n.'���O2�ʀ��9�s�7��sX-�q��� v�5'V�	g+o:xj�	5�!8��q&���X킖jJyL�p<�E/�-���Ȣ��b��b�e������^�B7�d
�Y��
�W�h�(��b�f��5��%X��O�!3�1L �S	�ܓ�p��Q@[���{55p�,�6�	�FV����aks���mi@g�����c�LWT�g�ҥ��������/M@��j���>s�������)��5�7���|T����! S��Z��K���m��[��ZS���������Fv��+6 ����� ܰV �}��_?ƱR�幪b'n�Ɋik��{f���M�AϷ=��QES��:uÌ�s�A�H1s�F�<���VX�����D�O����-����z�q|^r�kD0�"�@��C<��d7�Z����}z^� ��%�h�1� e�/����U�w�g{�>ꬡ�l���v�>9G����Q�ƹP�s�<�n�C�1R ��>��G�y�:I%N�;L!��5�rj���^t�YO�~����~�ʛ(�8���|A�w�ߥuV5T@��̤��Q�->`��K��w�"�U�o2�E+2*o�ۑgdU�F�  H;�"Jt`���d��̰�gQ��������#'3&���IAx7��H�����4�����8.W���?���>���)��M�eS/T�r~��e���4Mt���"hm��w���͆� ���Y�#��� a�keI��gʻ	��A{�!��	O�sPHj8���1c����j`aP!~#lc:U �h�Ġ��Ҹ�K���i�&�}cH	
��9d�e��Fп�����v��F�u��G��D]���:����
t�LY��u��ǂ�C�W	"�k��ռ�����8����Է��)ƕ�(C-ט>����+y�8Ins�c!�{�*s�3뇛�E?bK'��,�b�4�5Ƭ.�B���^�x�ű�U�bz��6L?#�;��;� "�#֓��(�/j��Rߨ�>ޓ
���S��{��
�.�_����m��h"]tT9��g�=��u&)�N�n��3��[ �t�&s�/����QK≀�`� ��֦gE 7=�5C��㜸�\�R���l�gƦ� =�h�U�%�8�_;��@�����p�;}e�ÊXcw�$H�)3kf�!T�hG�J�&��Zp�/gRNo+�)�h2C�Мk��D|cG�G5�|9v⁲�*�#6K�/��I8�p����a*���V�dw +����
��; ���	� �̾��_e�v�]=���5��'��=U�e�V�(�|�@c��e�<����@��?	�Oϩ�{��U��:5/�j�c�NFE�5X�#�ա��K����v4�,�29�~ZpF�+.Ee�M��@��q��ҁ�~��\��'�.��lP�H�˃�[� ��=���*2/��m6�ޞ�,���*5P����rb��\h�q�5�r�έ�~V���CW����N�y3[��ǣa�-Ǭ'��I��խ���2^W�A��� �1��<���&O��)#�\�g��9�ګX���'�P�:sn���o���k�9���B�*IЛ�L}V�W��/gj�3�6Ȕ���gR���10)�O��_��ܧ����#)>"�X�es�r��s��w�u @7��_�"������џV�΀�5�%���V"�% �+�&��rͽIA61\O�n�w����:�O�6.48Uk����<�k�Y.�	�R�L�#Ƣ�e�}#PGU��_��b~5k��LU�*}�0�tդ�m�˻���I��Y��-�o�caOj. � }ƣw�j�ꤽ�``SH�s���g�笾���'H� �ޡ�c���f�9�d�T��������@�)������لZ����,~�7$@o`�F�7ѭ�0�$��� s�'�5�M�ߘ}B50��Ȣ��y=Rh�3�n�RX�zdunW睚E��ܠ��ฤ��8��۸����[�@�v�3]�US�]�;������:�ź֯�=�uX��T��8/�a�2���)@��X�j�)�v7O���!�$!��lµ,(����p6��-7ZkȦb��O����Z?-Z �t��sn��h!]6��L�N �����7���J�G�-�K�0���Q_O��/�'ÀQ"j��wyi�?s���"��FX�[��5�4rˌ��������v0��D�{��t����rb�������K.
&�����-����/���g־�Z���h�>��HX��4`��?���1*�}"�!��ƴ*������33��R����Nt0rp+.����$�,��o�'F�>x���K��~��p��q%��-��bLn����*,E��&`�#yD�!�ѳ�������'9)0��Մ�]�pz�'dQJ��EǷ���`��`�{���&�Q`�֮n�V�>�)�W8��̌w�Ax]*�#h�Z�W^�3���II{BU�	�s������e����l�W��u�&��r)��MhQP�_�z��=��#G� �� �D7�ږ����%+��R/�<��s�jFJ@%G7)T�f�\��n�Ӈ�g�#�O"������D.��ѡM���PD]�W���5�s1�dT�����4{y*�Mc��$-C�Y'�[s�%���5��h�G�;g�J�(��v_(E�4�}M<y��g`��r]\���;m"�P_�+l����ݯ��>_ڴv3�v�'�@��Ԑc�q�s�grFw�I��!�0��*A!"3��@	�ӏm��*���� �#�#�?2�r��^�b(�%�gU7aV�T�Y�9߰/7̔�1���a��˥�/��1L�2��s_�2�2�/cqO�|�+j��{LU�Z�Bi���^+�v��Lc�E�䖛����BA�4�tyH���W'AN�2�-E	H��ٌ�{���/e�_�Q�G�o�gB���s���Uj�Dm,�W��я�7ܜш�N��}�G+�$G�UHb�����Y�'�װB�B���Y�N ����> ��YT�l6���O.^���z��,%�@k�%���Zt�_;6.���>r����!-u��\="s����C�3��-1�3��i�4"|�)�!K�-��v@�Ri����N�Z��n��n�� �%�2�h2�7$o��NZ.��0�i'����r4$�v���I�v��&�/���(�f[��e�`�����rQ�"O8�q�KZ,!Y�ܱz!9�Y�@?>^��}�iӁ��N�L:17T�mB�Q���*W1�W�ñ�^񎃇@UA1�D�$���
��E�e�>ī�Z��U��,B,˽I.ˑ�F��J���>��`�ߏ�;��?�̕���v�A�C�i����븍"�h�����H@\����R�q$�t�Z1�t��[!l���*�g�FOs��F��r/4���|z��/�߰{�Q��,�g�?&�׿Ho���)Gd�K���໎p�莎�K�&*�Lks�ٖj��F������ń �&�+�����:�J�a�*&����&e�y�f��h��rvR1�=���IQv�4+Du���<j��UZ�DGC�b�#��8��3S!��?y�Ã71*���=����kw4���"$�H�1������K�w
.]��	��)|��7�LLu��H |��6��a��"�fs�(P�b Ծ±�d�`JY�F�gO!/O���w�U�7T(;���o(�?6�3��Ӟ�f��LsB=��|�a���h�ӄ
�r�v�����jTO�+~��ͼ�-��"h�$�-{�E�2ݹ��}�x��!�_�5b.�陴ơ�OF�2y�^�`�"�E�������>O�P9�iv�P7����u�+K����{��i��J_��q3����:����+�ǲq���=QA��ݕ����=00w���0�8���#�{W��x|
GRMy'�c���6�>,�����I�K�K�Y���ؘO#ZbeJ��z���Rrs�)z��~(��C�;4�1;� ����c�=���2B˰�W��1��'c%:�H���Ÿ�:N��n�^�A]�+ݗM&�Ɔ�S�5S����H���fv�f��`�u�!�%u唾Ӿ%St��@����u�+���Kw�'HGN�V
���0`���¬5�I��3nz�#�\��ťxj�7�um�����(2����N����і��z4���干�%U�Չ����@�?�F��+���)��0r��6���N�G��!�k���Ȥ�����1U��Ƙ=����!'��s�F:�*��E9T�wٰ�������! �/q(�"�D����vz,[�B�L{�۝�6��J���a��GMl�n����v�W���E��[q�'UJ�Z����@0�&�-<K)2/���,��6'�=�4�O��Ք�Yݞi>~t9q�
9����|���[�x�Lh��3��cW��߿T ��U��hAT�J�G��r��9n]����bȑ����KNp�tU�k�I�*+�:��Uh�q׳%��9�p��k	wi֛��B����;����z�lU�*B�9�r=���=��KoEPI����Er�K���"	�lq���̀�I�.A.�F�}f���֍� �g��
�p3^Xqi���1�q���H�][�������m��-8�8��g#��|s�'�xN"�=YL���6��
� 2��/jk�l[]���&E���Mw�۞uH)����������	�-�O���Ĕ9��U�ㆠ�՟~S(�m��.�
{���W40�x��at���������wժ�(���N�����
x���O���Hx�����{٩��~�LjLR���0Q3dX0˻�x�[/a����B��$�>�t�V�T8�I�W;�IZ�P� �I;�}�j44Ta|����z:�#�W֛wɑqU�,1�����W��)���&�t����/Ys�����8�K��'(xX5Oc{�ubǛ�� 顼�.R3\�t>�w<@H:/�pQ��7�95k�H�=�I�|�fh���i�^WV}B�Set��n�M��;{l��c�C��
<�}�_���ig�訥�V��wf�O�m}��G��*�{���LD�@#����E&ozd��M��Y$D����[,�v$ϫ[�eq������ <w��c^��`�?Wwƥ}���|,�ԓ�?}��Ve_�����p�����ϧ>r\G�@H�r�S�^4VJ��i�$`�īv��P|��7�@V7*:�5��KD�e��3�ʷ��>-I�X��8;q�F��A]����#�Ύ$�[�2�����@��8
2g�0�6� O�1��xM%�8�r"ȿS�����dt����)H^d��n[(H -��XJ�>`�Ys�ţ���T�IR.��n�y���k�=�'��`��j�=�4�w�N|��/f���tC���V�g���Ȼ���M�"�R9�Bvnfj\FE�L��wO!��6��*XH�,�0/By�� �H�mV���;��g���1*��#��Z�Ɵ]repV�x���Hh��|���$#;�W"=�c� �*/���a�x�H�z>�q����=�O�ꞑ+J	������l��Y��RW (��c2dl�E[�GH�z�	djo�M$ ����{�d.'bt�T�## e.��J��Mt�}�.���{�y}&>�d�y��PI�r9� ����W_	���N����Sҳ1�*�37�lZ��3��-¡��Ob3�] �oF�̛�o�a)�����`m�R8�K?���I�$:$���iò���͂Q۠R����n��;s
�=xO�9�<���}BҸ�I����xzwA��d����Ȍw���ܾ��$�&N.s��K���Tu�����r��d
�э~#�5�j%$��>���1��a3k��o�-+*C�U3�\�+�A���70���(���u��U�T����fR�X�@" ���/�H<4A�$*�9�e����/i�a��##x��3��V�@��f��wF�������_@�H�����o����F}|(��|��.�YA�6��>�t}���qp9���9�]�g�X�&�i���=����\� 
@;*u��`�2��_����s��vf�Y�m�B!*��fe$���m*�Jp��q<:��0���9�;���)��[�<M���.Kݲ��[���;�&�j<ɸ ����I� �ϧ��s���~�
�J�l�W�l�eTH�6
>�k��� ��}��<�JE6z,�wZq�	�ӫבX���{�Z9���)-"@�"����Q�`b��'AԨ����?�XD@۫$TȀ����v2�����n�V2p�Z��t1�+�H�gMH:�5��>��mpi���a��9��iiD�q���w-�~2׶�;^{ɐ��Vv�IW��*:"z̳˕�;�&h3�?F6�{c�֝C�F���G��B#�V�CtD2�ܘ>�"$�% ����D�~�Ԟ+/钺/�aL2�[/���;��v�L� /'D�:L�oؼL���ӡ)��9�BJ-,T�,���&k��S˝�!�Xs�c�ƈ���r%Q�؉c8\�Oa!m�J����V�*��;�yU������A�nc lU�OCIń*7'8�kH����4X�tǦ�f=�
6��v"�r��P�k��U��W�f�V�W�y����&���X�<�(���BJ���U&%1!��y<A!��$d-���>�l�byܪ���;��,$���DӾ��$�[i�c��K�T�qy��(T=�c)}�x�K�ʂ�>�}M��+_YEjZ)�:M��>y��Y5q���Tx�U{Y�������[�L�<��{����囈Cr��q���s�]i|F�R��9�o`���#Cp��+�;���-���U����)���N3?B:�^�W��Y\������~Vrg۽��|
3i�A����Lǻ�j�E�ݜ�=�n��f����4�C(|P!Sd�~�ܛt��/����o�vjD,�b�N]�1;��=uo{ �<�+�D�:Ci?1����u��Ŝ��e�l���q�}���Y�,4l	J�*�Ʒ�1<B �Wjʨ!e�f�t�UV7ة���-��V��7}�~��WG�tٿ�|,���S�+��_�`�ϿЋ�(��3�)�ʝPk#�h�G�I,qVU
	f��$�:C���C�w��	�,�r��N�=�A!*�/h"]}:���Qg�&�s����`b
���~-������P����e�-+\M���Վ�|dLe�lq�f����E���'������K0�J�'V��i���*ģ�kt/��Ρ}��ׁd�0��`�'Im�ƣp)��e��ְg,�}��+ܡ)���3�t�|�%��}̮��(<���k�<AF�����(_�<G><�k W��+���E_vPZ���-i¾^��+���a�sm&�� �Y��rp�16]��lԭL3����<�-�^ROODq��4̓[��
e��b��������'r!b+��������� QB���2#��o��DW�H�瘅�	7���zP���T�}�H��@g�@c�OcS��2́�.�o�:�����s�5QLqd}j*s��β�Gg�Lo�F�Q�w���N��Y�R�II`_�\ڸc۩kmDD!�vC�:˂�v�e�}b9
��ߵ�� G��2���=��=��˄���N�DAQ4�]Vܺ1ԗC�P�J��))ͳ�$��0�1
��2���m@���G��0����f���[S�vY]N��HQ�4H���^�w�a�kP{Xf��6m�����!�ON�?)���-�o��䝓�s���A��U�h�B\H"J�����yD�S��`&w�)��l��oz�7��21kݽ���A�ݻ5��V/���}~�d��/�wF�r=ei.Ԯ+l��w���s�Lolxɭ�PY�-:?�f�H����=I��;���2�9o�/;�L�����E�_p$��?�'�}��v����@	�'�x�H����c��Ҵ>n�(�),�Y��ҷ�F�N86!z��q���A*�����w��7�E�dF���E2��]���E�#bb9Ӏ6���\��U����fVP4�E(��[�A?��fH\q(��]շ�����3j�PG���lt�Kg��h�[�<�}[ŵ8��P�)��?X�_!6��MEx�G��z�$QIb���8�j�i!�Ugl"O�@����JOH}=�v[�XRG�5aN�|��4d"d(m���Ņ��מ$c�1	�P�?�[nt��qi~aT"�ц(o��pӆ�H�>�Wt1����x	7��e�>�O���ρ ��B2�