XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��Plc"_��x�ҼhgBv���������H�YWG[4��c���J{�]_I�����x��� }�����G���F������h�xF�;���(���ₔ>G\�Ք�9�{~KxrA��T3���6�DJhH�$F�/2�Qex>��/��aF�!�΁��I��^/vz׀�gҵ��i�p�}st.��+�գ��|�(C���o��;���G�5ĨՉ	�}����ʵ�T�qL^N%�D���q>{
�]t��-���a��;�����4q�x]�G��U=8�lA��/����q������Y��%�0cz�����k�����T��oss�p���M��ϞCz�j��D Y%��ⷸ%���
\��v>�V>��{��>�Pm�y���2�J�� �!�V@]͓��f����L�����ǎ�5l�(˰o_�_���4�8��4������C��7���"�Д�6�m�Y=��YNݤU��}w[Y�ӒqauGZ-~s�RV��2IP�ҡ3&�E�}�4NU]�@S��[��U����Eޟ%U�\G�&�u*��������L]Q�³8�17�a���eB�f����`�W���)��.ڡ-�P� ������o�j�:9{���F�t@��A�?�V�T?�����׳RuG�貆�	�{�="G�N?
�|~��"��Y%	Ϲ���-&��/��k�	�}�-19&V�C�Z]��>��E:��Z�4k�.asLO�uJ	#�Z�/XlxVHYEB    9852    1d10a�#�E����� %{|���λ���fE�/����V����>8�m|
�1�u��?iײ]A@�D'����>���ۈX�w��~~���ėכ�7@���F�P�]p���/�; �i[�Ʋ��]�_H�xQi/O������b�bo�s��T�yG0�}N��E5�ލ|�ݘN\m�cr��4�X�v�({	s��kǕ��7_����p��ĵn9�,]O�;D���8��.Ӳ|�Z-c���GǦ*6ad�?�ie{�'D��Ɩ����=����#�HLUN=���3S�TV��G��T���jHܕ��_w��`�����Xin��8�Z��JC��I�{
2t���`�����9rE9S#%�����Ɍ��P��Fl�+�xH�f%�o�?S�J����H�N��ƪ�ӯAr؇��1�~>�sH�a~C�.R����op���w&����?�D��w��ɼ(��C���Rt���pgCyn�aE�>�����xKo���~�r3�ȕ����-��G6�������$}o�(u���0�}ѝD��K��V��"H}�X��e���,�r�&G�z��l&%��aF�)�l�j�$N�mu���S�E;����"����=@,F5�+��o�eD=3�ǉ���=�?�M���m#�-V�� �j������j���%���{@�蹙�`UQ�A�!;T���\W֣�Ñ�p�~q���� ��Jj����߬�bl
�i���D��YG���8v�x}C�Ayrtks��t�>dq^| ������B^H�zY��-�?)5Rh�}�u1�*x��U�ZFr̈���;=寀|}F�'s�G���D�P�tn��ʌA�5g��.��������<D{A�T߀`{������W�v�,��/e�Ca2avd�v��!t�ľ��m�}�]����~+WG0�A̹b��'���0�kC��_PוDT��fx�Hc_j����u�s����m���f?�cJ7���tV��J^u�X�>e��ͮ�n)�t��p	R-%
�����t�E��Ö�Qa���gdy�B�G�`���T�_�g�tX�?���T��>AgP�|^q."��Z��oJ��O��'�oF:E$p�:*#���}�mg37��������gJ�d8qZ��)�nn�j푇�/5O랮�ْ"����ȵz��\��tSl�(�bV�Τb˞4wB�b?�/��9��b�P��E���.�[0����s�2]T�����CI�+�-n=6�d�ҝ�h�� �<��7!�
���_�y��Q���X/��o�f�uVo�BI��ټ�`���� ��;������m%�nň4�� (X^s�}�y�Ef�4�O�m6mX��v�E���$+���٫h�O�[by�Б)h"�(����a��C�rp�KUY��\�E�H��
f��%�6���%���R�O�����)�ٕ$J��i�q��Y�ۼt�<�m�kI��q����g��&U��S!���Ս�Sc��zel��,���j�K9��!�wŒ��0,F�j�t/��io�0-z�� �
]|(�IM� f�Ϯ
;VДס9d�BW���o�xD�\Zh_�L7$N�+�+�>O����Z[�M���r����/�UZ��D;�	����M̃Э�����A�b:�Y��+��Q�dL�ܮߩ7��[�m�(�e/��+0����ʟ%��+ۘ�+m�*[�c��,n�sϵ�x�^�^����S&C�3X�~l�`��Uن�]-�4?#.$O=t�Ζ#Lc���O�M��waE�W�E���\�	��`k;߅��[��&� oI"*����4�����]|^U=kR)(��O�����e�o��+��0�m�K��+��Q�Α��m��7�aL��@8宬]�9�j��Z�&���X�.C���}]݁PAћ2�s�����x!g�`���c{�L�H$nD�h�6�����w�0$A�R
��{{n�Z5r�~�<X�un �&ȴ��ta���I�!.�E�8�E���&�Y<;���g,�u�+��8>����H)*���b��7�$�Ҝ+�-E�����m<����οB����@�Xa)�S�7WO�2R��#ΰ�x���ሓ��g&��D;W|8�EWV����#������S|%�Z�a0�#��v}��~�_���K&�׶� �Xd��QpbV�yR�#=$�V��=�h؏��Wd�5ɠ�T��������ϋ���z�2�ƨ�#2�d�H$��+$�쩕�j�k�v_�vF��U?>��c�ᆘ��G��	WK����i��Z��|���3�e�B3��T�Ry�L-J�U���A��4_������X���9�=:���8(��@����B?�k��aD�+��1F�h[��f�������c���,�J�����jq��� O�5�GVV���� ,P�10f'�]9?��'pģ&��'6~	PV̗$(�/�W1�f�����e%��
�"Mŷy@Y�in�[�1�/��U�ٜ,qV�^�~h��ȩ�)���=���mª�ĒZ'�i�����	��I���÷�yb6��wdVr�^Aʢ��/��N����E�,����T<Yjl�W�$Z�,^dk&4?ϳw��/�O�t�`�yt������P	׷k����&�,�ϛ|�G���07����tmC�xP_��MI��yh>�� y0/�ݪ�暹������E���5۱��H ���|� ͽݵ����>�4���aW�g�2n	q�:O�٘�� �D�	�j�� �[�d(|��n�
��Uk�C�L�iIe�nY�Uƶ�ǻڔ�LQ-���3m�4N��:�|Oa�"K�,zp��q�Oz2'�����/��g���m{����I��1s����"�'���b{�Y�jkK�X��^��,�Z����^��XA!��mo�`��*��5����.���B�e��*&�*��M�op`}�����K�A��L�O�E6p]���`�g��2�nN��+	yo���B���Ľ:e�Q۟6�2v�+��Պ��w5�^k�q��,��:tNa�J����z�v��VՅ���v���%L���z�c!U�Lzgq�����LrB8�����8�d�$���ݭMѳ��L���]�i�G��2M<c��2n��\~�P�.k���X��`"�/Ϭĕ�N|a0��5�;�Vڍ�hb�ɪg0�
�5#U�^�xŤ�9���^@VP��-��"JW�%T�eو�<�q��_�"\a��b��>I4U�[� O��)���@º��y��..7��k��;�&�NWqH�u�$=�#�^f��*���18����@��`ʶ�R�_�^kd0� E��N���6������)��nw�p��b���5��P���'����>}����.���̀O�J&���v��|���%x@W��4wm����	�#ef�@���\���eLs)����ށJS�*<�4�~u�yC�s6�0c|Q�.��R@��s�92�Pyxrd�>���h#%�}�|�cjsM�����^���B�["��:@���&�#�D-1��@����J<d6��E���A+2�j�����)�@uX�oY�$vˤ%�H��J0Z�=czIAM�d
?��~��h��Ă��91����Nl�V_5G@nPR���<Ч_�ZwH��k@x]�h�e"^lw8�	��=1@i�^� ��0��O0�H{�Q���ĸ�Y����b��W�G`�&�`�ْk�[�d� Fc�-?�Z$=�`��U��E}^�/?�W�@���Ļ�נ���q$�%�dB�;��4JC&�ʶ�;f_4��u��'�74q��(1�F���Eي(��{�ټ^�Ǯ��/5g	�CojtV���R�+rx�S�V0~�Mǥ�o��Ru�)R�

��++?�����!��A�N^o,����,S:���n���`֊~~����&��b}��+G_�8���@���y�>��f��E��1a_0{���L{�g�j��!�5oc�Y	��_�l9W��l(##�R��$潚9���:j�� ���<���ʊ�йYWE�'��ρG�Jc8\�{	�~�I�ꚀX8�ɔ#�*�E8���ò;����X�^6x�V�h^~��f�x��Q����Y�ZT�?�?q��Ǜ2�r����U�����0�Շl��$���"���c<�R%f���Q��g�}�!K+�'ù���ڕa��Y�(��Y`��
�N�[�nG��ϝA���H�K������J�E�=H㓵���V���R
��uYXϏD��|(VՃ�;��� �-vYKh��g���
( �"~Ef�c����w*%ؾi+ק�ϒ���ց�P��=XBT�˻dŀ@e��tO�Bw柞�M���e-/j��T�0�P3��Z5��2��s|�$*���N��c4Sɒ��4� �B^Gȼ�Kj��	o����wR�I��|}��z�+3��A��������C�"&'���Qk�n.:�S\=��B�ݥvۈ\W�=�������겘��hbs����vb����X��j@p?��"���@�1wFD%e�Gpԧ�
M�㨫�I8p��h_�8�]�����1)mrD�,�����:R�R������	ܧ�m���1ĳv$�^�5ţFa�1cS/C����T;`��JT�؋����C��t���#�֌�[ZL���RΨn�Z��5�Gg���>A�(�^ԕ�`�IQY�Q��=kE�M_�Q������n�֕�hpB��ڰ�݇�&7��g"�!����oBz+@���
t͖�|3\�0*G��}Fu|t�ü<����M��q��;���Sz�]~LA ���#�'�����k'���?��v��/��?�M��`4XHa8|҆ģ�_'u��J�<
-��Ȋ��d��TZ�#���QeНC哗1�]sV���5�hv�\H���3<������b��è����/j��(�_4)�cy��g𢽜���-黮�"��ԍ�Y7�P�b��"��Z7�ש�G�����q��e��g dh��<��Q�O�s��q�E�+L)�*�E���*��T�J��*+���t����P�ͯ�7���0���N������v����:U�`��>-ɝ%�?�����XC]:%�3���h�j�~M���>���A�#C'k�d+�w0���<=îvv������>�*�T��H��1� `SrQ���~s����(��_�������4��)��ʢ�6���X�1B��g��F"㍸K<�Q����]KE��#��6y	a�Q2����Z &�L��`SbHNE��h!h�r'X�&��Xj��[��� ɕ$YB+U+�֟(�7�պ`&%���b�K�
l�4�N%1�5�D���HBp,�(��6�� �wh��+D<7[w�*�� �Й�Qǉ�;��4@�*�z��9X��y�fQ:Ԑ)�>�v'Dd��{����Lq[db�$Ct���^\�%
>�����d���54�r��P7
��`�0��ޥ�B�1� �dp(�m�+8X6\��"�Qp��EWU���a�ƢΞ�7�ř�M�)t����+�^�!��˅<-e�cn� 2s֠,�U�$S�4�@y�ڼ@t�=~�xܽ)x�ܼ����ڋ������J�wA�p6�z���k{�vG�)Q�~<tkt4�6��3e`V������ȓ����u#�$�_$�tsή(���Ąs!'7�����FSv��&�P?�g�L�I�����5�pEF�����AT)`��&�"M���hAj����)Es,�pf��o�p:]ͼnA��+{�$E�J����j~��'��k�V$|g；yuh?��7���s���r@����|�+�s��Jj-'mri����-ҡ:���n����r�.$�4�^N���Ll��)�\ 6Ȟ�}��G���WޛI��IC�Z�t�ҥ1"�ă���r�����a��{ �*���nH��ޞ=9�\��H����|���rs��*���Ezt�ب�����:"g	>��Z��;������E��9�B�z`tk�O
�H�$�
BL�a�E��W�f��V��H�q�)@����(�&���P�P����V2�,b0�zNx��W�I�� j#�
~'�4�nj�7i�s�R�\���'�����f:/�����U6	�I^�o`"ՍI,�т�ȣ��B��
�|��hկ\�j���?��c5� z��q��]��N�Pry�yB,	�s�|��G��e#'�x_���؆���w�дfW�ܴټ�ۈ�����7?a5�_�2Y]�J$�s���ڤ�(s��3�\4�<��?n�[��%6���Ob��ж��y�P��n��s=�&���7��3_�ȥa,�q�
k�s�x� "�D�c�Ni��S���[B�ek�xY���Q ӟ�sz6��v2p���Cp_�l�Y���h��0A�q�A�e(K��}���ͤ���9Vl�ޤ.LD�[2�5DD��|�Vܕ������	
K�K��� P�6�cx���2��C�#cX��Y�yފE¢|��}k�}�y'a:�h�o�@�Zĺ��5_ gz|�Qy~� :�B��˂�7������R$�Q���Mb#�@����L;��)���Y~R����0�������������5��X�6��������Rw*z��쭕G�S�8k�Iv&_�:	��.l '̪nY'�9.t���P�7�"�'���O��ye�F��u(�C�N�}\��
(��wel����ę���.�{�+T��MX��W
�W��/�����;�R��7�`V�y<�J���.���}\9���ߘ<�5e��R����������?s��Lch��U6�RFՃTL(Z
��|��0���k%>��-l��b� �u� Sm��Ͳ��^By�����~gD�%5��B_�I&��ۦ�0�d�A���(����L>|��@�Y/��J!!b� c�su�R헀;�c=�F���B��M�3U�`_�c����֬�?��8�d>
�tjz�+�3�FT=/3M������K��Go1�x<���~Dx�f�w2}����]h�w���6�R�*"�k�IO��#Z��<~���J��'��$v�!��L�U��o�,��H?�ױ��B�d�,��_�i>��q(V�����cnz;���$4cT��;Ն����a� Q�����|R�M���G0,�u��dɛxIr�5Hi>�_ʤ��2p�_���C��=ɶ�#�_�v�d{#��s�r�}�,4_
��a�;ӳt��K\�"@�B�