XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��oXT����Z��9�/�/G(D��s(p+�m�/�{h�Шd�2zZj�2V�x��%�o�r,��y}ێ�E����.y~L����г��7o�p��U���㸢a�e&�:H������cn2^%	u̲%�����!�����ea�K%o�ffD2DKB��(ںPs�]�Oʫ�=)��<W��V����{C�6)�7�ȫY��Ў�.�R|P�\ʭ�*�|��^d���dǾ�g���^�T��r'��{�$�2��껓�,�C�]�vLM�#T�(G�7(�́�VSI�5]������<�1�;��D��{�l�S�u��w1�&�ȳ���Q��@Yʤ���Sz�5��,MPlB�b���B��rG���O u�S�R�5�R9-S'^8v��Z�&2�o��V�o褥 X ��(������A�(�����W⹁˜0�Z��&+=�oQ���0b]�MP���_6=at�C�pK�P!,a�3(o�M7�R\V���	 �y�B� #�s��?6Η�Z�fT� p��q��4�zna��փչ�^����C�m��=���}$�ny" �'߻{���*p0:,C��:�m�06�0�����CKr�HДh����#���xB�.���Da���6P��߈���a�5��|�-aq����sw���q���7���+��V��y�߮���R2��>���ʏ;�.!�,�vInq�DC<���\d�kI�2�
�B�������-�{��f���	Ї�{;�Q���C[�XlxVHYEB    c804    1960��0D�a�;if ׾�l6�
�:T�4Ey��:}/������C�ˡ�k�0����ʡ���\��5m~GC:��TRJ�S�o��Lf?J���4n�+ر'2�C��T�QEg���)s9@��!����H�a�==���W�+*R����%�^���B�� 
���J���ܝ.���ބ�U��oe�$IA���Q�N�ː}�n9�k�0��&��2�#����q#��:�?</��'�_ՙ���T��zW�WJ�SU&}GUvQ���CQ���ڏ&��K���PT��ǝx�Q�Pm�R�4�Mءs�99��;\eIX���R��~�S9T�.�JU�����_��fL�uh��m%��q#U*��\��$�f��J�a]�uy��K<ף�Ң���Ӓ�|�2S�X�i�?���Dޥ��D���IS�.�\�c0����=�����.m��Y?z��)]U#�����)JMv��9�=/���*�~*���Qy���ʞC���Od��U~gx�r>قÙ���6N(��]�K7�w��`h�1���4fGM=��gn��=�z]��8�C��H��+�-p~��i�q��m��*�X(��޲�tj�-Vg�0КbnG�G��ܦ�LD���^�݄��&7��x�G$˖Ī�Ι���>P�1Yy��`�,2������rÏ�<�.3sܨi=@�br�N}ʱ��|]�It<l j���V�;�׫�+����k�?�� 㡕^Ĉ�3�iv��k���CC��]��a^:O���=3�h$�Sͽ���ȳz݄�:�i��m�r����S�Rn/�p0�T��pөiۃ��Ƶ+t4���Ot#���<���W����9b-�C
g�(g�q�]��/�� ��b���181lS��I�����t���zy�;��M+#U#w�{f�ˢ,Uar�����*J >X���B8\�������!�qȍ�'Ó fe�!�[�'��g9ke��D�>��/�(��<��Τ@���+n�_�	����j�;�Mt�8���U_�Fń�ibaXG}XX-��������~+�+�g�T����~�:HY�Ri��%�!��\w�:��^�,n����>D�,�٧x�+�7�G\_�kY�D>�|Z�������F�(���<��`=,Q*�d@���ȪVQx�c��U�Ә/��Q�
��#�Cܿ�>_L�y�zn?-CJ��0�I��l𝪒�DQ ܦ�k�Z1s>[h�0�hr���ITSǚ���E��z�e|ӽ�ޏ���9V����ܳ|ux���̚#�;�E�44��H��D���@�
5?^��g���b�2��e�|��?�Ha4��R�c4�jK�󎔂��$�,
�Y�n#A���(���M,^7��;Ϲ���=i�oD�����0K$�;�{2d�Z�@Q�DfNmZ�q;�����*z����v��,���DAM��ix>Ԏ\W:rѿ�XrP��	�Fa<���@��"|�Dg�?,45
�[ �j���s�E�X�p��h�HzΌH� ¶��h�/�a2�_D{\o��}�K?x��P^uM��۪�3.c��կϽ�v�H�̖�d�+�}�Y7_��L��GX���ڔ;{<�'q��h��$׮P׈0P0�	�WZ9��Y��2gq��({��Lw�s���=ϴ�4BĊ���j�ow���^�k`��
˱�R�c��h�j<����k��%s�K���%�����t�x	�Uh">��$t]0���N�$'؞]!i�®���s;��"�dv8��Eu��u�w
��a���5��&^
m$��PF���ܼ��V��?V�h�YM�P2㓭��R�t9�ޑ(1nw�މ����k�P��PE����2���_�M�Υ�xM�.�Lhb��ZgÔԇ���a� � �H_��q ��.D�x�>��3�6�J���a bܰT]��G�ڧ�"	&������OL�4Fjmj��9MFOKk���ջZ�$鲰������g���Z��!Kgq��#�qI�"�p=o�Qz�vZ�P�Lэ���1W�w����ф�/}���ڭ��+�RF
��{����l�@�+��J������
P�2�ӑ�Z�>��!J1H�KB�۳��ټ����b��9��{g��X�c5W�ʡvʇ�SS+��ǒ3\��B��x�R��0��bP���y�7����@C�i�.7�g����	�jZ*5T�]Es�#΍E^<d+A_�b����u�ȫ��9-G���������x�S����,o³��6���^�l��C�:�Pw<ڴfu炂�3�&���_NMp@��9���֣7�
�@�?Jmօ�>��~	qT���j~���W;6������Xk�D;��A:���Y�ɹFA`Ǥ]���ΗE�a����9\����;��s�ٞ ��Js��� Q����w�-��8�� �Y�^6�|����s/���2�	�n��}�{��m����齹T��f���'�@H���~Q�Æ������և�zx���<����g;��ɹtP�z��^r���f	�t�`˻�xE��;�Ȃ6�*Id[ �Y'^wl��꾶����-ӕg����(|p���3������;a��s�ąҬv��[��$ë�M&�(��~�������zk����z�j"a=V�_!��g��-i�qZ�+��������y���V���ߓ�����{|y�V��&S��=��:?��u��![�|X�Q�Һ�=���m��С9����
�g=�gR�D(M:R߾��e{Q�T�����X��jM�{j�t����gj��>�	(r�#���m��jee��\�c�0�U�M�ɤ�=�C@b(2I")��_w	]V&Ỵo�%.6EEOra*�[CC
`˫�Z�Rm�>^��q�����赩��Ty/�l��/����"06>�#���\a�O�2hD%k޶�B�X���LH)�XߴwI\��A	�% *U�T���b��K�,��������T�>�5�l�?���xX�1�*,SY?�VJv�V��+}�E����e��N;U��֚���a3��6�#챑+SA^7��Ey�� �g�0�t�6�tt 5wWO�Ƒ��Q�G];�tcD&�)��ߪ�!6�PT%�ٜ݃���+��h�򘟴�5�c= [=T��1�0QgrV���/���U�{]���N@��A�j��%	:��XhK�	��q�c����I]���~����^�z��5p����Η��&�JwR��N	��ɱ��R�j��n��f��]���A�bNNF�@�Ѡ���niap-���_��i��!�zR�(:����>�X����Xy"�-�����VgfَW�Jkw���ݶH���J�ޮI��t�'f9&�v����:��K���,�ĝ#���A���g���z#2���x*I�(�,C�<do��U��:RV�i���նA���Bj=��A���Ol�َ��fĒώCi�@�L�ϛZ�(9������a=���Q+Th��U�;�{h�L3���?!j��8�a����3ݍ�M�WBl���ǋH��I���`½�S�1���:�WD0|����|��^���Q�]~�H �G��/ۖ�W���V^7>�u+�|��Cp��xI�����[�-YY~�EҤ\��	�?�������R�F��؅��t%�������Ӓ9d��������5fp��IB��su0W����֞K8��geI���^Ctu�!���
���94qL�W�@�t}fx52���>2Z-�^<����͊�կ��n������w��ye�X����K4p��vF'�ܵ�+���;��Z�B�U�&������3fkߴ�:w
��8,CĜ,I�#����%����W^	�?��7S� *P��a�H�!&L�ҭ�~����7��b_����sgN��/CE��M�D=���6�	�:�2{�Ir�d�r�P���|�^6�\wu���}��Ǡrq�pN���y�����^N9,��y4W��R�[�u&�F���k�{Z�\�{�ZT�L������am���^�"��3҃Z��D]��r xT%��2��+�t>9��_^���NJv������Q��6��$������hP:n�#!};"����Z��[��B �+B�lb%�w��}%�%�F_��cO;"qb����)AdP�5x�B�t�b]��.S�gV7D^VM����X�\ڹ��"�V�����S�ٱ�t��� �#N��'åsh�f�g�Ң��Dl�;b��V�����U!�y!h&O<�Dzs���DE�1��*�O����`^e1v|c��3N�ҩ�gk����"�u (�vʳ����|+4x�7�6�����������>=)��5A9t�5#����#�t��b�\U��2[.X�^��#G�C(�?�[��,m�֪�p�o�q���R���Xx���\�����H.u<�F�Ѭ������Ů�#��|�6�1d�hW��Q������q �]d~�pjI�Iܷ臉�S�3x|!<d����UsD�V�<X�b���$�Ί}�yn��\�`D��*�&�e������O3�0�����\�cԭ'Zj�I�Z�ɶ�
�5��ZS�Ǝ`��C�b�5S���:�-�l��SS��86�Bu�\3%�j�iT�l?i�]C#��*��H�ǚ�=����z��p�x4S������佬��k�gl�s:X���}y��j��۰h��cdF�,
�(ZTʚ���U���st�_Jg'���ޑ����)n�C ���#��8Ί�su�#V.#(�p��/}�T$�����om%�	@僽���R�S:�vE�2	S��8�49�ޛ���(Fɖ�*�,���6h�A�w�z���4�t �.�p�~�?����0=Sw��F�r�گ���V����>�� ��Q�9�����H��жhr�(��h���ӆ�*�	�����,�K�73s3���9�`Hi����U���7O����җ�m��M�Ù�e\��b�0�1Gt]  ��\�8��C=MBX0��0�/�ޡv�pd�!�)H��.�����`����H?eO����<����'�\%�lom�0��;R�L�N��Κ�xg��$?Yp,��gWgr��H�S�-��Ș����ҽ���T�RZ~�$��;z`�6�i��4i��W��@���x�=��c�~���A��s����kd4��Tϙs�����c�_ýo����<n?�z�4�~�1]w�����z>�Ƥp���Bۼ��{�Vq�����dC-�cF��y;w��/��qk�K����,͔*��!���>p=o���e+O)m��\S��!<���ux�x9ەeS���e/$���jSқ$,�GS�Gld�DrhM��_j'�������Mr������k+nn�ɽ^F��lO�p+k1��i{>�8D��K�6PI�"J�ܭ�m쎚J�b��wU�d7K�.�aK��K�`����l^U(m�u�]�J������Ij��r�� wS6+ӂ��Ͷ��`�	�����P�v;���o	<�i���L?�%b�X��Xŷ�k�3�X@���<y������Ó�|Hc�����6ݟ�K��u��/�nXf�`�9}b?<��l9���W��
03m>�Dn��B���t{~��'Dm�7������(gn��>z�I)�������%���6Dt"!#J(��O�1ͅ�]Ĉ. ��Һ�Z	����+�w	3
7G�Uj |��:הX5��91���q3>�6<K�9[�n�\<��e"E���{��^<S��͕1�
FD���;�F�u;��Ϥ�v�w��A��ɹCa���9�P�{��Y��9��1ǗK.�|�G�s�Ja��q�m�~����ɰ�4�G�ɝy߿�q.�&A���^�#!�����@�u�־-�#<�}Q鲁D����Nϥb�U�y&�2;���61��&�M����A`7��S#;B���^����@�M�ۡ�����=%���g�p�� Sz��$gꮴX�2�/�kV FZ�wJ �r-Xk �-h�z���q^+��ndvl��LD��>R'1P.%�Ӌ��\L:���ҷٳt� o�ȂY;/�ז�Q� Up�ÃV��.�n��M��������=�W�@�uy��4ۊjao1�?ڲWv����Z���x|NZr �����-��N����	��裐1�G�-j��"�ܞ�ȶ#^��ք"!�:��E����q+�f��j�/@��(��s���d�Q5�D�IƣH�Vg=����"���� 'D_Z�1����ZvyE#��qNC۾(���͇��tôN�p2�������<]q�ȤG2t�a�W-���