XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���6�C�0ta�s�wɒq�2@�;9i��@���ɚ�4�(,��\S۰%w��1�����S�Qh������2r�Ӻ:85!4Jm���%҉�V�*��q�N����g���16M �Œ�G���Rb(
�KǊn��Θ�u��rY���/no{��;���/�蹺�)s��bY��a�Ӕ���;�����b)�����g�*�8^�x�ݐ��iD����5�,�������>7�G�W-W���3�^��H��&��8�)\���=}.�.r���@ K� ��b��D)b֪�;V;���D!�^'�k�wT��#⌡6p���W��rb`_KG݇w��^���x���2�Ľw|����8�C�^�ŀz���i_j��NqJu�n��ܯʞ�����V逻o�޺�Mw�sEh��.�9V�r�M�������v�����F2�y�%�uj!*�O���@,0H���1�E+ށ��zY^�;���C��g��B��O��ܑ4ߐ���8�u�B��oY�5�|Y���+ɐ�����}�Q�l��q �p0�4���R
������$~8�XBW�e#�,���;|�����&�� `#�������s�4W'�<� ��a@��";Syȶ��H6�|�}��Sm�:z��,��Q�-|�FN10ݹ@�/7�]�X,��U�g$������G�L��sz�wJT�{Q��eW�X*}Mw �������;$�o��=��j��XlxVHYEB    4284    1110�,�����xt�`=�(��b�s�uuR�'���DB|i����Ak,�� l�`璴���	�g�� 3��P>s�4p�N(�@�HJ^��}8
3�`"�ר�L~x�Uޓ��W��xQu�W��"���<��#".V¹�F�M�Xf��l#����]�Zj��P	PթQo��ͪD�^e�	�+���1T1&!%4���T�� []>�$��*�}[� A8c�<��b��<���:v�z��B���p�~��)���&���Wc�cCmǊ�D�������Ϲ���.��ϵ{6���_�1O(�4���M���-t�`	��_sʩ�`/G>�dRP�>V�.M�]5��o��$.���l�"����E�H�%!����л$��Z�tXR����3���bZ�Æn��V:$�)w�x���Xz �TU���m��1����K �ȋ�%ÀE�����y=�H���ͷ�$&���N`����U'�[���2��S�NAZ*3��U�m�1�62۩r�I@�&K�V��������i���vh#�t@��_U;��v)*$��IIі)�k�ˌ`ЗQw�V�(U�]�Cґ2l���-�s��ނȋ�9��c�R
��$����w/j��*����N<��:�,�.{a���Jo�3�w'�o��;��/m��\��]>�2? S*bi�I(_�`E�I뇤�]�3A6b����-n�Frhc�n'��)a���9�1�\��)m��-%&�9�*����$i�l���C)S��X£^�	�[��F��lB�d�������}Z5jF�/�pՖ�	��1lM"���8���# C�K�cԠ�UeQ�́�q�QB�p8�M�����GԀ�At(iv��My�$؊S;���BQE�:���I���,&X2��B�vvQ/��D�ֈ�q:f^�A	�I�R���T��qUp�I'ɸ�b�Ѭ1�{�{�C�r�p�?AՈϾk�`��Γ���,��,�N��{���4�U���)�g��HY<#6k�N�B|���Z�bz�Px�8��o��x�Ē����`I8��k>q^C`-�Oo���u�����C��%Xk�!:>�,ǝ���[I̙�.�������� +^nz�XdL��v�ay�C��
:�\N����R81RYؙb�B�5Ξ*�b=r�#�W04�1��dI[ƚ��8G���q&F6!8�=�D��N�����m�d����%}���;�����]�,����8@/r��h��E��ΰ��J�<C>C�+Ω� ��!*i1�ŏ}Y|F�p��e�`��#����̳Q�A���<j1A�<��ȁim)��/���y��)��S�!,��B��A%S��1��[\�
�8�鏶_�Ok�ϊiXx,�ߘj�-7��n�&�-�����_u�P���~�t�5�>���{)4mf��3��(F:��{�� |����F��EbI*3���{��Q���\�v���G���gbFi�����r{m�̩���9���k�j�&�!R���xk����JM��s��N��e�3�Y�cw35�yh܁��x��	؝�0'V���.;�Kz�bOk���r��d;����Ÿ%E;v0&�ۺ-aŀD��E�#1��8�(-c�rT���&'n����_ķ&�~�:�m�y��U�-3sgZ���K���)�iGogV�(^|���Z@�k���V=�	Q@�PF�$�֢���q�LӋ�D���|$��s����ԁt}�H7�ǰJ��E�r--�n|�1J��_*��r��M�ߚ`{�0�+T��E���׎�"�c#��ʼay�X�AR74�����,?S�Kds����9"Q�/ݻ��r7�\^�Ajn�	b1���nE`�,9%���ߌ��x�H����m{2�6z��xҖ�_���#{^�7���^����ж������5Lk&
��~ �+?G�A[U@	#0��(Ma�я3`-8ܮ����G���Yg�ڶc9X���K����@�}�)���\6�*j8��ϛP�/�Ex�\�͖��L�ު�,�L95�A籗���w�$~���Xz���⺵��NSVD{��X6.�D��h[R����^!GF���W�0Vbwc�Z����_�R�5�J�?���������D@��u�2s)����׮�����ޑ_M]a�~X���!d��`3���3��˼��+֥�#5M\8�Á�Plܢ)'f��r.(�e�yo����<2c����/�f���v&�~�:��Smjl�y��^��ΧCw;4_NAȀ�4(�v���"hp](�h 
�.c�e��nC�Q��EN'de�����d��>J�z8�k���P�L�2 �� �]k90ֻRv[LI�����ǂ i` ��e��F�Z)`�P��(�$;&�m6 7X
=��Uq��S^�Qr#�*�S��k���-l-c��a:HVa]\x�G���}����`�=`QSo}T�P������'�s�c�kF�7��)#n?x�<E~D��Ɇ�`*��5-����N�=�Ծ~�w:�Z�}D8b��<� �5�Dz~ԟ DS��o+OA�'$R�CG��l�AM�VG� �K�~�.-lT�Y�+2�'&��7�vסK�RWx˗P�9�@�/:Q��Y�d�P�6d}0J�rJ$�i�-��m�;�4B�*o��Ҹ�a��"��m��V�lZ���X��3�*Bb*ئ�i�ɲA��-����Q�K"?�c�{a]�ε3OÑң^����n��lr������*���*j(Rw�����э]3Ѯ{����J�q��Phs��C�[����ܔa�;C�|2/�Pq��j���?_�[�W8��H,E���<*���0N���>�x�XG�����l��� _�:S{��F�pbhh�'��&/U0ŕS��kDB+�
��r5+`>K�/��8Sz�t��1�>�n_Vx_j���d6�dE�bw�sJ��pq#���7�I�ɆGZW%��̕�׎A��P���+sN���\���4DC8��g�嵉��Z����#���)US�K�ˁ���|MN�m�!����rAw�y�a���$J��k�n��ǔ�Vcm�]l�uC5�	j" )�� Md]����#�Q�~Od
��v`?V�q幭���c�v�����.�։��`�j��LIJJ�|�	������|��@��I�Dk�nH����ф5F�u����,kS�l�re����SS��C )�d4'$�<襲��̠U�j�k�s��و��[�Nȕ�8��	¹��R�'���NYx|9�?5N�ͩH�R�7�*��M��6%��0�
!��#0��n6�0@#����"��9��:%�`��ܑ�{�<��d𭏂x�0s.�>@f7�|����T6��# zs
��ƥ+)I"0%@+Mt
U����Z�Z�X��c��u��˱K���8(��uҷ�Ma_����;Pa_���������7���OʓD&}����#�~�~��k+�N��~�ŋ�.P-�k�SI(GJ#�/Ò��W�i\�\\�S�z�S����KUW���Ҁ��)~ǖ�S�-�h�9�
2��'��5W�e(���<<��z� nI���
!U*��?`y}�s�):��'HmR��.��}h�掳���
RĢ�Qb��[����1����K�������!:�{W�g����d����-�	�^� (�,r�Ce�)3f'�U��|��g��kA֣����}e�揇��Ѳ�pQ[�a�Pc�����y��h�A�1v#zǼ��ul�������yb���o��aƵ�<9w�e���A�W:n��{��5�ډg�ě����Ǒ�/~c5�����L�L'%���A�X9�J�c���>��ET*j3�r�Z�b�A/2MO�����G���	�=*jj:��c���jC5B�I���x��"��ӡ3�s��G	��qĦ*�q�B3r.=f_��F�>��:O�L�pf��[�䀴ѨO�X%7̕�/�{����V�>��|ط�� 8�DM}�L~b��?�T���s�pמ%�ҟM�������v��a�׊�.�6�Ij0�PzA�d��%�J���{����Y�_�/����s�:�f��xp}����~��(�wv�{��֜P81����%{-n�����7D��i�8`>~n=� ��i�*���"����l�/2W�1�������UDI����6�ly�e�Rh�MÆ�	*V���!��!sv��Bbx_�p���ជ�Y�m���B�!��b�i�|