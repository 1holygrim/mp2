XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����'��Fn7B�C�Jb� ��`���fО3a��-]
9Pf$У��% �5�F�#�`�X�ųk3dw�SWڱ�/��:F۳}r�P�|0�E���!3|��<�}���|�p���e����L"w0L�r#\�p�>$�*n|
g�$�"�	Gv�Ͼr��UD��\�K�Х5%@S�D�ݧ��*!v�KL����]za�ϳ�ԣ,�Yڞ��*���q�L�q��v0��ۤ�	� κ*D�aG�w#�H���(��K�|(����^p�f$��e�S��Cӑ���:�(x4��H��s���5h��0gږ�Z�PO:Ҧ�9�.���'|����څS��g�6�dil�~�U�@EH��?C��%d����'���-^;��69�̀1:ǀ����~���,#��ye0ھF'�x���ys��&@r��d]Ek����x�>LD6ty�X�CT����ޛ��^Y[#��8}��ʀi�����%�հŻT��� ���'�i��	,Ĩ��w-N��\�#��!�'~ր�<��ea��Z��S-�E��c�eD�Иn��`�u��)��ѫ$4�j8�-f%��ɯ?%\+�l_�t�0�n���2�@��ޅ0�U=��\��%92�ն����O5J��7~&n:����D �#u�]��̢����ɝ �s3��4C�BHG��@ 
n�EaW��Յ���W�}�4���^D��S�A�x���ϞL�;Xi���;k��|������>΍�D\ܥc(i,IXlxVHYEB    5224    1740 t��c��9�����۰3 >�e�ZdD�=֟-\܁�F@p�]�0�R�P�Myn�������/�kC=ӵ���&��]_�a3&�}�=74	Iɺ���ZK`��[B�4��3�o#}����F��D0B���V&�r�?���կ9�C�O�7��c�%�"{��[�@�h�%[�֪���boÆ0����AnG�nۊ�у�3��{aC�/�%��(	���}O}ﭦT_�:�i�p_����=W+abg�%t�$�yg?J:�O�_�N�m�1�V�&��D�;����f�r_�%�;頡�'�=�݇:}uP�進��s�H&� �|́�����m��	�p2�9��5�H�֪�|1��(N�y^O�*�Yc��۷A �S	[.��p�<�����s���оʁ�1op��yj������������0X�~ZA���j��D�\܋hb�.o��/,�t�i���lF�	5,E܏V��z�"#���~\��VJ~��(3��}�!��h�!Mw��b�w�V���Hi������ޔ�w��v��?m���P�R�p�3�܅1Q��fm=��f��" �9O8.C���.��-�-��D}xR��=��3�	z�[v_��82���%FI���])573~`i��{3i�H��"�����.����Ǚ�0��W���#��5��Y�`�);��Zm�-R��(�M %��U?7�㵪��}�� �iyEl
p�+��ܻ�D��2�GJ�g�T�z	��%�M!��u	tSʖY��g�6�U���[FФ�6(�^��dTȉٹtЇ�ЉW`�J��Pn�%���Z��K}h���8�iT� �pQP�&��,��P-[;���*l����Ȕ^s
����	��B���oM �Uօ��0��X}%���TD.|������Zx�; �@R��Wn̹|��uR�l��R_���`�&�~��Y��M
�v�����#�AE��k��W�?F�$�6�߭D\�N��xE�oR�XQ-���9�;�:��av��C�G�Y�����&��� ��TC�i3^:��B1��㩒�G믒1p��6\���JX��Ã)�r�	sǒN��oQ��j��m}c��D^�:ƻB㶽&�-b(b���T�PC�e{��;Ag�ˮ�$��Ìw&Y��vG"�btD�&Ð�%��p�*SZADbii?����&��<�%]Mg�pm��ѣ��ݾKS�B#���������(��r%P�cg�c��_�w���!,�䟕×�P#������MyZ�f̺h���Ѱ�ob1��6�֍K0��R�W�#�c�	�e^P��]��?�a�%T���������}���W�9kj��0��zZ�%ɪ�(_E�:<����jG�ɭ�nb�쓎NYV�Kv�92�lt�/��Zr �e�RƏ���*0̢�i�����0��0������v�����B�#��K�{���hky#v|��)g�N���2���a��^�]0H�G��h(
+֞�k%�^bO/�:���`����
|ћ���c�qW�}�+j��Z�Lhpl�I{@����
=&��?�~�3����#	�0�v)3��dʙ0X3�u��L$N�̀��r�EeLJy,og�%�?�IW���p��E� �E`�֤m�۔����6\�1���b������e�]z���k[�q�L�6^�Ɲ�?9(�G��0�9k �z��2.�|�nǮ�l�IAi-\�~�w޶0�.�/L���=bg��ỻ���ah"$ ���\��'1@g�-s$"#��7����LQ� �zo�CŶ�������Tj��Կ��dP����g<���%JYNn���F>r�k�u��rS�����_�:���3���p�	!q�)��{��z˿���컊�R,�	�u�"��1�Z�Ƈ�T6mgN�����L9P�h��׮��
���O �<d�x(���1���n�pP�Pf��Y�2M�~�ֽ$*��Nw�h�8
ŵ�h.Q��Ը�!��Z˒���v�`����2���A>�N��>;�[�9�!��t�,&�u�z��J�E2��꼇�T`&E�\,�1���|!�����/�h�����R! ��[8�~䡶s�\��S�K�!���[7�Wa�Iϧ�r]�x��;�mRGC��,U������T�v�Xj��Ү����/&���z��oKҎ���4�}w�����Y*�{b��B:�<r���z+��$��$�fuP��m�JR���C$�߈�/.�D�(R��bo��d�|�l+vɔLn��'��
�6�$Y�*v�05���K�����Z�4J�4�m�T�r:�b�Da��#9��<��yT$q}��pt��	��:�y=��� �Өw����G�Q��Э����-�Q��F����|�\���:� �R�<�B�/Z�vWъ��
�8v3˞�Z��g1H���ْ�.S#y�O ��-��6��J�(¡~Eٸ����A�j��J�o��*��ud���"@Kr:F���=d�6>2��H���`d�_V��l�jEw,�A��U�z����5T�H��f!�/I����wN�U0��^�l9]=YIX�R��n��ױ�wꩡ{���ju��g�q2.���?y�&K�Ĥ)���� ;F��fc'�E���6\�q�̲�1ls��(�=aa�v�npI�S����!y,f)�9����M��:�|T}f���(�h�}���@��.Z���Ͱ$F7�u;�:��IQR��%8sKQs��P��$q�(�ή�n��%�!G8���VDE"v���_#����".P�5�A�j"��)��&*�Ur0Gv���<�X��}��	�?�1�Nq���$�x#P1:?��p|�BP��{���II��;���W��ݑ�������zN ��Xվ�R&Cк8swvU�@�`���#�M;��Ԅ���/�j&.�{zА6\<4L�����c9w'�|�K;�t�J y;E�פ ��#�����=$�F蜤Ux!nTb/�X%/�J�j/ 
���̉u���γ�Ԥ?�z�)�oy����ld�cη�zȉ?�͏HΎ����;�����bK>��v��<u��s�)��G� n��j�?P"/�A}���.�X+9��ð��},R[�o�@�����x#nQ`�ifR��ڽM]�1�!&�Z��!��xp�q�0-~wc0�������o�)�s����8W�V��]�8�ȼq�� xV6�U�#��5��������^��׏)TC.0�.�;�\�[�~�4�݀�{ QO���^'R�,���<h{��n�_��`U��/������a]L�
U&�LX&�:��E	�˾4��C�*����F����Nr�t�_T[4y'2]�j��ڒ���8�Z��U��bF�j�����x�(��r�%�y���:ŭ�x�R]�?�E�	��p�]�$h����Ul�ؑ~�I6!�I��a�o�^�'ǆQп�/���X1:�ʖe�d�Z�B�Up<�?o�^�ې��R�2:�ic�h^���TE������--8R�dL�g��(�p�p ���8ڟ=)d���]��c�EAB��<<�+o��<�yr;�T$X�Z�C��x�?0�p�%@�V��
��t�ѪAl-��J���B�Y��-�M`���\^��]���o��/�b_���>0���Q��S\ ��ҋ�z��ȝh�/���J, �F�` g)N���R�����;���ܧ->��w�t�C�©��3�V�ͅ��Xw��G���٧�g�!ĄA���o/|e�n]��������	V��A=Ҭ��_X�S�����z�|�G�`K�&�X�u��T +N�t!�b�L��|�F��#	��L|M�s�z:6G�ɩ�AM��R9�8)�m$��n)'��@�Z�#4q$�t"�ZM��џUp�Oj5)V�p��|'N-,~Ot�K���L�g�R��i��J{�K���@�酷�\��>QY�V�,��t����UKa �՛���8i�#�k�g�¤D��د<�跅��zS�;8�ݤ��m-�%��e��������T�#��H̥�Ĝ�9�E��`̺n�dt�"�� ���S��|��݅��H��S<�7��Ų��=���꤁�]mN��i�K�Dʰ���e���,�k�8��׍v��v��^DA�d�D�Kr��XL�q�4�M$Hd������ $��j���X&�*_hzN皅���y=-�Q�̑p��K�H�	R�B�7�u=Y$�>�K�C.���vN����8����C��c��k�>vd��p�a�� ꭩ%\��(�*�/sDw�/��Xߟ��KD����q��+_|�
�L��2�:�QU^z�����X�6��Tː�T�0IF��*Z_���m���F�s�$�����5�+���:���o_h6G/��h�/e#՘���H�8}���"Im�K8<��lt��z92-�F�O���F�fz������v����'�녡���w��i��Xe��t�#J�f��@�|}-��߈�*�P��^��]癱>*�5�_�Ź2@��lI�Fm�/N���tB^��]����,Zi )���]�K]k�>��G^p�he���y��(�y�1A�$:7*(Hh��J�T@�?��e%UH�i���O�8�P]��D��D��S� �+~Re��r�x�?�XE��[�d��RgoJHr�#-So.�h �ho��mo�c�ט�� b^<8�i}o�ɤK�+�$�Ct�p2��֓\Wr8�V�j�{���#����� �r�Eʙ���(���u+j����:�W���ij5�CN$��`6}O��_.Y�.�HsΣ[���O��
8�Me5���i�'[e���yN��Oi?D���:E��k1�̊�l������ p��Qq)7'�|!�")���viF@[JIV܉��DFcS�kHN�?I���������93}Ry���=`8�%Ǘ���}�`\��R`��9�(�>��Y���)1�İ��e9�	��P��k���d%W�}����b��+�Ԕqy���"w���/s]�/k�P��0�`��i�>Ճ��{W�g�a�� Ih�,���g ��ra{sŰY[�����n���)`8���o
�!�C0�F�j�-2&�VO?�� ��[Ʀ~��o���=�z�䂊�4x��*
�ͤ=HI"�c��o&�PI1ߡ�d��%���y������_�Ezƴr���;I`u��/V�5�)�b��p�⌤	�A�*M�拮1��!2���AK��<B�-ncv�;GEB�C�C5ai�'��.�p������K&��������ھ��/�5�,��x���Xg�Yaa�s���M^A����kU�h��rjɎZ~7	A,����V7���Ai}��vZ=Վ����P����>n7��Y! hLu7��i�OL��_�-�B\�l0�R�߼��q�u`MNq ����\P�6M5.�#Z�������
�lH��A���K���n��74n�0s�Y'������S(~l� 䘻�bPf�Re}���L|q.{�$KmQ�؎CI���h�Ub�n��O���
JI%x-��K�wRؙF�o*��:\N����v5�7u@jh_�,�4b�_N.��)]�^a�g���EW�oPI�,ŚH�)G҆��PI4(-f3�h�]�ܘr����R��ܺ�@N#0�2 ��<<��%N`�Em���L<I�� �P�� 9O��m�,:�I/�#v~!� �����g�>��F��@������<(�2���E�y�:��׊=%�	�嶄�u��m�z