XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��?vg��doA�/��(<B=+k�#�ǺK�jR��S1GU���
��k�䣻9(�VD�[��"��2Q�z��e�\ph�,@��C��hβZdi�r'��}�nd6�4���Z���ھ�ߥ�ߟo���˻dݖ�R�b�8����:�
c[ަ
��!0�Edg�1�����s�*BL>�9��^��H�c�F��7q6������]K���ׁ��]��B�A��޼���V?�xԹ�������>h�i�Q�?��[
�����!�.^��W��N�)�B1������yH���ˈ<!H?����A����{>'2��"5��W��%3��|��܂ϠH�񁺗MZfy]�����5�W�W�Ps1���9�{7��J.������Wa0�4b��g(V�~��h�}�ђ��b�9��z�j�B��z���+�T���*��FI��-6i_��lh	!�f,]���$�<�z��e��M�^U#|;�Ě���w3��AfZ���T����B>:���m�*��2�2�Y�x���w�9�1��n�hl��(��"�ٲ�&�8
���	A��8[��+-0�b��T�uIR/!��������a�|=���b\��I�#��Ͼ+��:T��'���41�����i�o1<ƴ�nF}�ޚB��'�U�#�A���N*2��}�L*��o�?���w]mb�!�~5?�xZ�s��n�[����;S��|x˾W�����sW���2u'��O,XlxVHYEB    1f41     990��Q�_�2ۡe��=W���0�k�EY��Ƌ�A7���n&�&�Hf�?�p��MWK}��b]�W
�~������j�������0b�����w�ӽJ^5o~�\�
�Y��ӥ����� �\�i@7L��k�ظ���LFj�>:15���?%Դ���ŀ�ֱsʓ��I�|�U�4�w�i�W��7D�{�#vs�I��hߌ�O�Iġ�r�1����.�^�����C� �$��\����:\B���P`
���Qd��P�c�଀$�qz��w:3����[�Y����S&���h�#�D���� �0��� ��1[D�\$�m���P����R�O����7V�=n6�?�����U��p�5E�%Ncٵ��4%n|�����N��F �f������[�vB��_�����ɹ]�=�}�F�!a��A\�IL��&���u��lݠ���T�8�d}*�����\�̓�O�>�uܹ>`����9^��x�E�1�5�h$��K�
��Q����_��(,[�+��؁��SJ&�ծ���#(�L|<���fS� ��Eȃ�����@Y�[�
p|��G�����e��e@�,���L��߼�ogQ TH�O�a�u��x���W�I^�1>4� �0K/�Dꬶd���[!��>m��R�J�E���da7MQtj�t!�K��Lp�\�U��j�-�.UeNHJ2>_-q�<}ne��.r����_]�q8��R�U NyԈ9�d��t��*��`���p�p�uh4���r4J\K��v{"�Z"�䇼 Q�ֽ]�dZ=
o��j>�EM
l������3ikh�p��x�n��Ѫ� ���1�?�:|m1xie�Q� �*#t��W�s��Y!/���a��J�8:���WoChh��CA��Dt���k�����I������I��Rݶ�;� Uk>�f��U�$�0w��.Tc�?qYd�^v��{�`Y[�Oe��yq�>_)��\�:4A�mtÑ��ɧR��Ƌ�g��5a0���d>:M�(���x}�jl}ʉ�,O���bRP��3Z]PѸN�.�`[��0	W� ���(e*DQ��J|3$O�-�TES!�� �~2g���4_`���/�b���a�qzx9Yi��L�Gm��/QGJoC���^�O�ON�	O�7	I<�{� �����h6s��	<�`)�9As��@LD
�Yy��-Ƃ��քe�Z�V�s��~�qf�ŭ����˓1X3"�S��B�J��D�-�~o��5�}�_��Z��(U-����4m����E��`5�
�T�_���o���ea��$�֑ԋ���tP�1����wl����,G-}?[��Ou���O�'�2�2��m1�#��y�||W�ti8& ��0�����|d�񉙱"�+�aT�y���֨��?S�����^6l��]ڸ����I�2��a��gXt��;0&D ����>��Q�� � �E�����ɳ�46��[&�1s��7�L Y%@l�G�<"A��������VL����,�d������>iG
���3]�WVK/	� ��-��W��i^�~��C��uuB��-L��e,,C��U\g���J9<�Wi�N)ϱ��������lB�6�/��$�7L�)!��R�>F�5$��C��������y
�n������E,$P�.�Z��dž��N�hٯ�w��ps�c�Q�62b�j�p�ѧ"��"�s�&���ڑ��_)���O�ygKY��)P+d��{^�#��f�_����f6�cR]
3��F9�9'[`�{;���>t���m�/��l�K�Tl�2h��7<���U�7! !��c୐�\ɵ�L~���~F��׽��7l�h�!b��Ɯ���F($]w�-�R��:>k�����؛�<�4����՗~X4s_qi�S̓9Э5J=NG�}q�Rf������F ��CAh�R�^�J�]�X%�ܻ6����:�m�{�EO��}�o�	
*����)����aW�[d}s¯!�P��6@��V���5?�h-\��Z0>ǝ'�}Ł2�h��8�h�\O����#�'�.`��\��_b�O#+���d��b����@a]�q�_TV ��hA�>����/����ӣ^����O����5�[��m�;=(�qo��:dp}�M���%��	��|�m����K� q�<�K�-���ɏ-9h��V�5�ث` �O�)K
��:�;�QP��m}���;Ҕ�K�4� ��Dc� ky�Y���V(�N�;��W֬?���V��������BV�ϒ~��G�>��+ @��=�QxN�nm�	PSNP��e<f�x�cj�;��{/���kt�f*���z�r�c��Zi�m�35e���X.���
c�%�q���܈��l0� -�