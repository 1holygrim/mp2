XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��Pk��蜩\������}���Vժ��TM[L�=�'�3ѕ/�LM)iǉ}w��L�k�fj<�ǀsi����K����pPoF���S>�x7"jŇ��fc0H��	F�ⴑk��`k�7xX<q�i����+:b&B �ra�)2A1�o���m�t�M�Y߹���k0��DS<�Zj��x-я?���^,�:�k2�-C���s��7�8+y�Eh�M�m�?n�G�j�G��ʹ��|�D���_�\��]�Wsm�՚0 ��e��,�㱉~zt>�S���X�,���/�Ԫ���~뮎3T!JT�:����ir�B�����
轞<3}IC}B@��/�/YL����d�'�ɯC�:ٲ:rv�	�(D~k. x�/���ؽ�˨^QL��w��%��T��087k����m���R^{�ߧ��"-M=Un-���r��x��Aj�p��B���(�brFp<D20�G�D_���)��{WüN�_����\	$ʲW#�B�w�o_	RS*�L����"ym�u0�XC�	G܃
�M�t~��l��2���Fg�����Q�̌Md��R��ߦ�E��s�3��@��D�8X�W+Õ|gx8a��Mv�QkEw����I}�}ot� ����d�\"�y<i۬]
��a���o�2iĀ��;����D}/b�>��4s�2t�ύ�.T~�o��ܢ���N�2�k1�jy�#�Ԥ�Hb��9��$�k�$
�R����>I���yP��w��j��XlxVHYEB    c05a    1dc0�@�Y|*ܣ�x��G��F�J�#c��M�®͉�ӵ�r��
����+9]X�[B$�R58'l�F��0�?�cj>U��36�?Y�hIu��q��'��)��q��q��Z�>o>)���,�l��Fwj��	p7e����ᰱ>�����:[�"x�*����d��E�-�#���y��] �y�Z�n\�-u%��ܥ_v����]bUKi�5hR�O���0���Q�$�6�h�z]��OAo�Q9Ȥ���[�)w��q`�%ۀIm�t�"�^���-�j��R�Ԃm��Q����羭P�+�����b%7�΂|�gͳ��鶪t�钄6�sm�T7��O�/td��U��4�q����E�!K+�������&��Պ�PCi��x�J���<�k�q�O4�O����E��`��׬ۦ�����bf��4�M|����5/3��"u�(��L(R�����[�X}D���o�T68j��n�1 �*���vi����'40ݰΚC�?�C�d�R*������1(Ӕ�NDx�
I�I�`I0�J<@��S��BTd��!7U5�ꔓ�g,J\��
�~^ǋ��e�5	�N
w�6f����b��>P�7�����~'Y��~-�1��ШW��x+H�U��L�����	�n.�͘���fLU���F����&QvC�g#eԒV��,�@�����7>pMc���ma:���]JweL��rcvo���N��'[kho�A(ۨ���'+G*�����tϼ�n�~P~���m��W !��D��WȐ���"wc��ҀhBCCa���,�L��;��8� �A�ZMv-
��>ۘ\��+�3`��K��c�OsZ���BG�F������BZ�w;�1U&��="5¯fE3ky�R,>}��ݖ�,!�j�]�f�x����*Z	s-`N�f3��)���G�����oy��]��C�%��r
|LgOK�]�������4F쬐��r*��\u�Hɝ	�����p�b�1N��oÆ�M�'crXD�(���Vm��_)�b�*��!ﴃ��P2�j�v������P�;���u�ۄ]�̟x�����D3���٧����_Zm���&#�f�:Z�(�Caĸ��9�CD4B�	~�ެLm��f��]��4�2��{AO�Zg�U�W���˙6+WD˷���E��dO��i�>�o�n���2T�7e0[�?�յ^�p`�Dۛ�ٴ����h�S@��5�:����p;%������X�lkj�:�$��$���&�DI���O�$���Ob�н&�F<B7����Vm�Y-����6����&���4���4� A��*�f�R�N���О�E����6�诸��Z��1{3�<k;��
�=�����@�i6���R/�2Qz-�?�:�G���.�,$��X�'*p =͢z����=��tW���Z�%E�}�7�<HP�`Ɩ��k��C�K@�Y�J���
]c�r�G�x�۠�����zbNxP �FE����Ǉ6�	��rU��(�a��$"'�,��s0�uʹ����i>�I�ȿVmR2��Kc�QE���zŰ.k��d���ϫ�c��'Lݍ��K`x`�~��-�S[2ݘ�v�ᡓ�3U�T�C�����1�5�c�����v/�v��(Q�
�e�������~꘳U�}-?y%���C�7�7G�~�"���j>��a�\]W��tp|3�h��0{�9�w�<Bm;<.�T�,g��V����/C��x�vW�͏�<=@*3�؊$tk~�� ���pH�8��t�A���������T�,I]|^�?X���̾s
�	�Nܤ��Si1���c!jri�$�ۄvf��VD�&�����;�bÕ�yU43N9H�@�q�����P�N��s4D;��I��G忦\�F�[D�@�ã�\�rI���|�!��&җ�HWl��	�˵g}��� öz�ENV��i�W�NAܲ�G�#u�'[^N;+:����rI������h��=V�OkF�GS��	��X�y��i��݋l��8c.�U��!=U�/
I_:�i�AW�}0VH[.�S�n4ؽ(���Ə���k)��}ީh"p�^]I��Loe��خǅ���ќ#�?J��+*u�2~k����|g�6��8~�g�n��9y0
M!��(h���nn�v�]v<���C��DH��a�N%�}���/H	e�0�p`z]��x��TU��~X��@�b�SJ,awo
�<�v��+�^�.���^ׂ�z64d��n\���R�k�/��V�|�{�D��I
=���3@�)��0v@2\f��tsyQJ���/�:�<*��JO�����T��ȑ��G�З;ۘQX���5���.������l<���P��������O�|���J�im����鄳Y�~��C����� ⾺��_E<��"ׇ݁�?��~Q��!�7��sѳh�T�ʛ��&(����h��o���>74wwe�U�uKtMa�mHR���x��8�J�nQdh�1�9����1��RB����}qg�D8�[ɿ����DFqO��y��{���\���
,%.g�f(m�j)�m}qZ`l/G�ߌτ�##�=Sz?��� J��I���1�~���ٟ=�O~�E�[��|_
Έ+�}�Bf��x�R���@�?�?dmiJ��PWV�o�O·��&U!g��T��A����_:`�K���<r�%��q�A�(�;	�y�*����C�؈,㸶��5Ӡx.T��!I�"ƺdu����-�/4�p.���}�G�ߛ̴�������d���6��?S�|X��Ink� X�d~�YB�����t0�<7�@�
h�ހN���39,0� W�R���������w�RgVdKζ�-6g�z�N-A�˙�'=��t�v(3��`�^���r�jPq)V1��H����^�]e�Y���cC�����K�A�G����&��2$"��!xx���;`fZ��H7'���U�oF�M�FȎ��Ⱥ~e�̫��eZ��F�_6�푮="в?��2$کԪ���IE�χ`�V���`��,�NX�)-�����|����,�1���>
�s1ת-��/���v�:�|2_�WX�늵� �B���y(ld����)��	��8�����1y��Z��6��B͟�IC��Ɗk�|��O��G�Ե�5Yn�bE�?��6�"���S�������Ѳ?��L�$��ձg	{B��[c�G���@*�_��*�2����u]��DCڈr�u���h
9�Ad]�댿���픸�_3
��W*6;u��oH��oX��v���{}Q+�8�Α$�M+%bl��~A�����5��#ʾQ7e���EO8D�mI<��s�Mxcjt�.���-��P)�n]��j)LQ��q/�9�=�PG���QVA�3�b��//�GERbKC
׌�E���69ũ�p��9��Y��CioʶZ�bC�8Q��ڨ���z��Z&����}o��\�ۘ�y�5�T�vI�we�mĐ��Df�^���[.y~FZ:ٯ&4]��J�]~������m�_�0ܓi���k�otZ�Y��j���l���|tzl�h�%�f�:y��s�x�Z���y�g�b�I ѧ�]�rHH����4���^��$�37���sQJ��ҶE?�0MS+�L:��>_v�����.vz3-*�*�^;�lRcP��A:��=��J��k�mǯ�d ��Ja�Gu$���R��w����}HJ��Qo�bg�K��|{gۥ,�y ��E�n�/4O���Ç?%�����`����[����s<�^ǵ������}�����YBqy~`�5�+�ʩ`�?̈��9pK!�2E�f�\�8ͳw��&��n�rA����;,�^w��Y��q{&����p�7q??Oʗ9kڋSa!���,�rT@*@�{4�j.'��8c�e�zkn���/��K{��0$c���c_=���*�W�=����0pC.���'��~��W�d�ߛ�D�i���ް���Q=}K�41I�����]�F��K����<R'6��֖�~�4:>N���J3r��rt���u&z�<[{��өB�4N1�&k�е_��V�)H\ 5�^�r���w�l�<�)�[�/�yA
Lt6�s��G��HN�����ȬE�$��`�	eQn��Ƴ��8�7���ҥv�LIb����d��M�ul�ry�,Yc8�����w�����'
��}������j�Է+V��(�e�N���Z��dy)4ઍ/��>�����~^�FS�>�������!�l���1���O���j�tݒ�9�3�}��7[�$)K��	s�$��>��фVII`.js��R����4�r�a�`Y�6N��6�2� �2��[U�Y��EQ����(�T���*�t�pE,S �Z�)'�g�%��\�%�#�G�����_� �D�AW����p̙�2��и2N���o8Wxh��̓�uu1�K{��!rH�o(�i�>|j1W��~f@��d 85�z:p�
��b��X�����<qnݛ�T�[˾�s��^��"�D-�<�gV.?�0�-Ya�B7i�RX��p�\�۱��s��zeiE����O�������7�#x�%yM>h�؍|T�[�\����a_��!�@z��m�.�s�t�p6݀��#�3)�2h%CK,�_���#��0t9��H fހ�*2����K���
�}Y'���'n�{R��S����֍!W�)ޙ@w:�<S�U�����nl�HYg�th~^�����;־��'����|x
�#0�s��ak�YoQ2z0o�^����+�1E2U��1�?�[v�N��p_��s�<h�݇94�W��ZG���r��7�3��ŌF�:$ }1�Wr�I��H�7J�͞PT����K�z�N{N2k& �Y��57a��[�PW�ЪL��јN�L��{@�-��ԱӊM�IT����Y�D��at#@^�H̡����Ow_��,����w����oR�e���~�&q�sq=(����s����1Vr��``�<=&�yƳL|�;d+a����_��T ��@9��X���8o|��d�i쀵\F��cmZ�$bF=���57L�H���-����,��� ά��K�*~�c����-=�r��.���Ʉ��%�3�`o�ʿ�o�0�.�����{֞�?�f�������S�,ٱw���:�?<�5�v��ۆ��łHI�l�_� �Z^�X��B�k��E=�=�1zS!�gs#��K�2���=Cŷ^����!�%�Ƨʘ���z�I�.�uU����#�F����w��l֓7��7����55�
����a��H陨��U�o�.:��A�
F��uڰ�]���TbಁQ���,<��z�|2+i	7H����r���H���R@�����yZ'��u做x{r�e)KΝyQ2�!���M�z�	`v��HQ�Uz%�4z�t�!�Oi�6mS���g+�F1�ٝ��ߗx���u�#.�j���K��q�?��:�ģ�$��l�,2C:]��b������J�iO̭���!,�bs�/Nc�:sP��&ޥ��0����:vC˔�elf�*�~�u�#�WU�^�7�1�����z:�Q>�ؓ�^Pt�i]�u�����x 8���A���j�vo�A��g㏗I�*G[�~a5��
U��F�<��	��q��?*Qj���S�T�-j��s�6�X1��Ji�:I����s
x���������kuWy��ʢ�AT]�(ɻ�=,�[]���4��KDJU�����W>_[�O���@buL�dG�8R������d�w���/��&Sr
���b��ʋ��*P��H��4��7_��E�e�J��k�4�0���ysJuegJ�,Z=?���c�e�y��\�E��F0�Y��:~��s�c OA�#c�hpwh$6~�`n����i�UK͸ºo��E���t���Q:��miK�k!�$�/��}5lUC���8����a����-'�f�)q�C���j�|:"��/�>d������j�N�Y�n=a�KK��)��I���ܕJ?���~�,�<�>��E�����Z�ؾ�{�e#��|Be:e�#�{N8���_�E �������&;q��fI߇;?���^�
��	�t�������������Čќ�.��$�9��L]�f�������8�u>���\�#�U��,���`�E%����6�#���V�R<@@̐K �M��v�Y�iR5F�}�u=y7V�'����ΞE�';����=�r�/3!�u�s�c:�$� ����	\ui�\3�"��+���x�7rZ�T~�{}qئ7�b]?�+:9� ;3�0*�=CE��-H����V�LLYR�6���E��|�=Ocv}~�/�hD���ք����;���)��]&��p/�3�Z�����MJ#��/��$�/4��A~JЯq[�s} ��`֐�6h�숉U.���D����q����Z�c�e@�6A���QJ� �H�D�9���������)g�\.r���+��c�:|��Â�Z����)uPOv-�Y�G�����T�� �+})�76�4�~B=]���$3�qx�rR�����2̒���٦(���J:�ކM5�n�VXo��?_�$���5���[���h=�9u�vZb��.
ZRA�Ju'�ْ$����U�����(��!pA��ܿ�6�]&n�<��Pj�6,�f�ِ�ifj;M�{\wUK�N�Te�#rgE�E�%-�̲{ ^�Zӹ���sy���#D@a�2�+��/��xm�v��� �%OǄVr��$��5ϱ�����"��f^�J�nߒ�����P�#/��\M��N/�'Q*�>d=S��������7wD۹v�����#��$u��k��'��<��a���Z�}�ldKk�s�Y>��4 i����O_57��h���eႏs'1
=o�i���uT���A۝��zd �)�u/kۚӪ��4\Z�ޠP�UK������)m��%��x��2R݆,"�u��Q�0�#p�x��r���>�+n��u9������G�,�7{��$p�??Pw�h��$��a
ے���o��ȟ��F��?ɯ�:�4�/me����CW-�M�^�Q6BQDӅ�&�<o�^�.�t��z)(�sV]����
h�����ѩ5�&��+���\�>���O�z�<��׶��k��3�oy�Z;�?����: ��<�}Y�n	El)�2nt�9(��U�0�wMޯN����p��+�y|zW�7q����zlE���9��y��э�Qo����ZJ��#V�@�^0+�,�F�qo�qCEhb˟�]iڞ�Ư��u��#����Кs�}��T�)k{�w�:J�F��e��A���؟��iq8��;�ޱ�=�ؙ��88