XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���I-�{~4�!&�>RD�@)��%��F�Ԥ�9�w��o?�
s���A'�}�mK�"���|��6A,�5��-�|�*d�����lm����p������ÚR�������<K#��� q��I�� �/p��Q�������	�����nx�^�W��2�%jGf�篜G�I>�-;��B(yˠ�"A�*��� ������?ϡ	fs��>Tۤd�I��e�K>TCϨ�
���������,!��#��N�ƾ���+�ќlc> %"��wwȮ�%�T�*�z@������v�-������ -��' E��zB�@�O���N$#b�r�5 ��/W������ .�+@�zz�����>��v�n_�EI#|t�W(O���C�؎����r�bD"����y�q��JN �s��yG�C��=�ǿ��f�[�%��Q�!T��!�:t�d�g�g���
� �z8��D��c+����d�XR��pX<C%�0�ab����z5��Un��1��ԅ�Gj���P�]n�Ok���6=Pd0��
���PM��3{U������B��-�^�߻��C���H��]oؕ~N�f�Y��+�S0�]rW	��U��a��YG#2�n׳����Áw��	��E��ȷ=�S��$�ڒ�<3��\+��s;ݪ�Ժ_pV�߲�b�����v��m�p*�DA���m�kl#�zEG%Nn%ϷK��VvU��Y�ј�^��c����"*�\�1jP:XlxVHYEB    2ece     b70s��Z�Lk!�I��\�\E;�}pAKx��|��p�g��&�4�$Ȗ�lf�z\���9*Oѫ�$E�pG
�bD�H����%*{�a����,9�sH�v����k���]>�1jB
�Jr�3'����(3��L��c�ǃ:��[��ͩˊ�
g"I��y)v�6cX��)�%2�:��/}{]�kQ�H�S��1s��n�S'4�
%:U��� 椀����T��[杹�pm��� ���Ў�#-*��>�����~"����[��~+l�ɚF!�8Ӫ �5��	��H%R[�aE;��������|9��ˢԂ`��d�������2�������^5I3�V����g���Y�u�hJ$J�B�Y��KCg3*�_ͅC�R�|��.�6���lI�i>�WDӹ�]��`N�����M΀�-:�7d����}.m��e,��~���H��	R��mو�Q��{n�fu_4��^]J����*�3X�;차حܩ���dG��g���uvQ��g��-ZG]ҵ������\ݴ�%݂��ZA�<_���ɱ���m�6���y$��.������3I(`I|St�'�Eig����'�S"������.�f��@Jv9�9�tv��'v����rs�)~���ֆ`dT(�hȹ��{H��$&bKk�:	�6=z�S�l�Z�hn��u��m<�#�Id�󉪙{�q-�@e,'R��]�x\8���`��]ޛK���vk�tL�v�B!������d��gQ�We;v�W�e�2G*�!;ۛB)�ND$|������3���N��<���c$y�uh���U�c��w��~��������u�M���<����/�bMYgl�cyY�M�K�7G�-K�[�%�)�oj+�~�v�E[؁�,F�bjW4�օX&{���	�#T���NM����Nw��k=N�	d����NY�U���{�p���LMw�\;�XO��zE����o[�R�ߊvɅ�y�,($X=���Ff-�0�{�]z��tٚ%P8�)�1c.�R�U,�#���m�Q_�.��N���w�rf��'Q,GE�Y�b���HDvf�!'rv�-@��Y0R��HL�#��b=��h�Y.<�1&|���Q�xA�����`�Ƕꜞ:JJ]>��~zp�\>m0��7�q����Ĕz	� H��ʦ�p�5]��L��sYT*�tS�H:�gZ��$����֍2�6?�����?���e���
V{�J%�F�Q�[����o��kg�pĂv����P���(,��R�Ҧ����,�!��JKM33[��6Rx穎�m�Lp��m��0�x��S��Q�mܫ�t�t�^[�C3�(�ݧ��΄�zQ���7�Q��_�_�&�����Q��� �H���~��rx����b3�������ޢ��8���K#�2�@�nbu>�giC��r�� �X|x������·~w���r8A2�+ނn�uˈ�|���7���ޢQ���*C�NR�2�kb��p�<��� `�+car�%X��s2]�Q8A�y/Qsz�mEdPr9DG�{i��Μ�@C_��ߡ�r��HZ�N �L�e.���<tI�ս�|���M� 9������J]b�X't%�=SQ �p�V~\�.{["�Y�
��vG����;'��5�$�M-+�?(�J���?7 Y�*|p#�@�)Ϡ�����$:�Hw1��[8��Hvo=�Ǧ/6j�ݐ]OZ]!��%W�"n�|AxrX�V���M���^o_N��Nm8-�n>�����K˶��"�����$�_����x:�)��m��Do��4�h
�1�ڪv�%qHR��?�5dZ�� $"miM-��2�����Z0ʰM,����$�n`e4k���.�2HI�W�֓P�Ӫ�w`\eD�Q_��ϙ4�v�ϓ)Զ?����|50�S����N�)�Cٳ��w� �I��Z�r�ֵ�%��};�R���d!�<O^}W)�Xt�v�h��B���r7C���ĄB�܇�*ZJ[�|��q���e���:�q����Z���~�;��9�+� 
�7����MH�� ��z�#����x�!�����c��`@�a�IIE��,�uAw��`�~�')�]�)�G
�8�?	j=^-n�m�MJy��$Y� �%L�5#��&q���]g��ܻv�.sw�S���F)־�	�w������U�"��9�q*��l	��x?�S�hW^��/F���g�U�y8��M�
�WlF5���oKu�O�����@�.��_k[5�2�2��� ���őHn�zZ�!e�8(��{l��sUz;ˈ�ܲ��Yq�M�7�i��R�Nޘ��� 8�H�zK��N���c�&��>����m�ѽ���7�Yq��Ӛ%��[�z��0��w�t?s��Zo����H��`KTJT-��m%&�Yifi�(���;P��a��k+��V��?��e/�'���]%���8�?? �{	4�_�K�ƏV�_��t6��KEX�$v�?��}b���R" ��'�t��X�$��Z�r���$�9���>x��5_���`�%m�r�ǂ��T���i�Q��Eh�d�E�)1f��c�0֗�A�V��B��U���a���e7�ן�\���%?��!Bj:��� ey�%���]I�+�uI�p�=��b�M�f����|��B��u�;`F�$_�H�x�tg�&�Y���g��Q t���{ʙ���Ϥ����KŨw) �E���a����RT�$ڔI^s�Z�*���$�R�oj)?�"��Y�b?=�h_�_B|rj�F-=i�A5���z��p5.��s�^�\�2����꥓�1Y��N���{J/R3�z�Q򖲾ԗ�=�*wP�