XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����ؖ6|�ثty�|X;��R �]��GΓ@�0�K!!Sd7'�X؂>LW=V�\^&��u��MS����ҕY����v��%�/��<�\.�d�Y ������NYon_Q����g��1��� )_���\T�}��2�4�U	�"&���xB�RS�%��^G�D����/����fH|�4���/U<��'�(������:d u=}<�Z��g��}�	��5�����t�`��܊#������?��BH�"X��C��\���Yp�q��j3��"��xJ��+��e�)�V�=T�aƔ�6+���G���NH]� ����ؙ�F�l��$�j��Ϟ�L��y��c�?SQ�FdC �$N����YӀ�Cu��wƤ�W�2V�v��s ��IS`P�����ƿ9��Y~Vy�i��e�U�C|�m�_m�U�����\ �VK��>��!���l}��rX̵q�K�������Ar1��j3g�y���1�(!`bD �����<85b����,r8���MY��MK��������\�G.`��掃�*�n��B��L�������l�'$������J���������d�:�2G���,s�0B1����@K�g���A���H3��� �;��ν�7 l�:�V�ތk�`Y��*Zd��Tw�^�[�p�٩)�0��?��hA��$BF�./���vt���l^q�`��o)r�Mrcr(	�2�x��$���CV�H����a����ZXlxVHYEB    5fea    1830}f�['�`D����.
YQ��d���ܨ��W}�� ;X�)&��e�йH�^��(��H)sۛ �y����<����W�Zvmi��C�-#ǧЊ��R��q�K�g�p3 ���8�h��zp��c?�t�� ���'L�����xcQ	�cl�o[�_��`_r�պ \*s1�]��3\�(��.�u������� V�T �Bz��8���)u�M�N���7)��:���8��A�ŔR/7��lQ�#��#�jU��t6�H?4&��^e�?�dƕ����;���
qA-��֚S���Sݮ�fyQ�
����ɰ��h�!�-�bpTD	�!��r���O�搪����j�2�V��Gx�
��둂��%��a�&��>j��<�*�-�z��*[M�>Fy���d�.j��n�>��C��2W�b���#?&�9lI]����1� ��)�QD+����kc���LW&����CE◧�?��9�x`��G(,0���cFԸ���~��iSr���2���nEW�]�L'�Oe��L95�QP�&y�e�Y+1�rS���͇1�ϗO��M���i���ٚ��4�E�x��A�ln��5K��4lg�Q5����$~a�w�W$��8-�>O�H��x���َ�{�V��>�%�_�\�#��+Κk�&�#��p
���P�̛���g��n�)L2�p��U���,)mX{@�Ͽ`Ui�)�3�����DӬD"�Q���[�]��oJr��7��!e�=��a���*����G�?v�
5����.�E�A��P:��ۼ1�My鰵ȓh;$�R��i�W	LQ�ӵ��B?0�L ^�%'�q���x�P����$�%\�o�@d!�J��8h�����'g�-ԺW�Ε��,�Jr�F��Xt+{Uܟ��HD��t�=���$�e��Z���*��Bt�+��q�2�uB'1���;�׍��b�tI#��+�kUC��ӶmyX)43�,�9�O�[+|�Ŭx0O�����2a�$�Z3��b��Â�t^"j)�^.��i��Eo�7�t� E�b.�����{w<�.�>��ۻ: �/��/���\O����	͝�F� ո�1��g����/�$�K�_#��S
�a��pޡ��s����-=N!XV���i�w��D�(�ٱ9�	?��t�b�K�H�א�,�.P�_5J���7�s���ls�t�s�sI�Nu�kT� w8=<�"0�4��-�jG�/��%�m��׮RZ�X�����<�a�G���#<.\D�`�7t�P��g{D�WX������a
�2���:h�d5��$�XpJ� �\�C.v��4Tz����$YƤN���3�U7��i,xz���^��}0��	���H�5cq��r����	��hm��"�xŵR��=��}�.��H�H�@HU����f�8I#W������'�= ����_��ޢ�y��M�	���&b ;�L��+�p=��}"��wp��g���"�%Ә^Z��x����q�N���n���
�zxGʇ0�9q	ؚ9/��L�	As�ׂ�Z�^!>M� z��w���l�x�d� ���AĊA$��h������4Χ�1<�;:�M���b�&���P��`�[6��W-�N�Rl���S)ػTK�P��ؚ�O�j{\j���`^v!�N�w�ˇ}��#��1��獌f斤&� �j�8��4���>���Ds<������`u��=ڮ5KR@�<-����Ύ/�����7�+L4���`� {?�|F�	���J6���h%.H���������(H�pz8\�yY����vv��n"����Ҫ���� k
�QrD�S��\��vmk��rhd��E�e�8)��Qp	�X8�����������Բ��m�U��n)n�Zu�\A��C�k�c�Һ
�/���is����f�,)�H��H4р-�E�t�E�/6V糹]7��r����W�oT����"C�y�~�����6�m69	1�;=ä��o���H�r��@��v�=cN��ӈE3�vE�ʏ��wp�<�H�ENa�0>���T^6V�;8�Bz�Gk����l3Վ1�r�7j�?�']D��.�a�<)'�NC�]pʇ��n���.��	.^���G�Ȥ��ɳ�4��i�>�/�u���aڶ�f[�洝y�%��,�aGg����*�hWrd*�;�ld��������L��s�َ:<�����G]�ض�6�8�"ó�XY5m3K�S��k��]#�ږ#���剷�#6�~�=�el�+�R��8�d4:}6��r�N
����NY�_��PJ��H�0�~՞�I|�.�ܠt�P$��(�]�^&2.z�Q��yEɐ��Dݥ����j-��������!S�0Yy�:�W�xk.jkN���T���	�%����$�v��K;S��G\��M̘&O|t�\�դ6'm��İ��}j��[N��.f��
�N�i������������@� �n�#l�}�縕`�Po�j�N߉&2��˳�cڎK�$\�h3>,��4�8�J"����o�O��
B���O�o�ta�r`�>�K���캗�Z��/|>[HwT
��6�3Q� �{���r�	t$��]t���"l���1b���٘�E�[z?s��\��~W�-�_� ���J�#*�P46ţ��yC���r�����<^2�
w���=אӣ\<�A�S_^
UK�N8|�Q��l��O���������O��F��O�����Wu['@��xp�E��f�2K�x>�r�<.��S����u���Tʥ	>�������Aw���o��Ә�a�}��^5q$y%�C�`ۗ~x��3����߮Ǒ�$)�+��oL�4��|u�8���>ͯQ�jp,I��%��������`���<[_���Z��_H�?k}Sޖ��T�_�������A��XF	�@��>��
�u������0X���i��$�yw��f��翉�T�D����7��M�f~*�3>���jD�;�V�n�߶f�Naui�	_v>n�9D���Y+e��<��g�1��3de*�r����Rv8@�V5;}1?�U�'e���#:F�i|��l��5Wmn�`���t��bY ��c*��A��ra?��yWǲ�pFn`����s�v�2�ek���s��8$$���$vf��J�^���c��c�z��zh�Z·�$�����D�����N�����&ua��BZ�gU�}��S�Fey|t�cڑ���b�����T��`wd=��f"���
ȷ�"���Pzfp1_�[Y����3��T�듔�3 t,�Tx�~qy|�p��4��٩���p'I�OI�O�6��~0�����DL6M� �������"
L���� �����ց�n��7 w�j��N3}mX^�G G%��nz}�� ��{���)��;,D�󆚎�R���,D8�[�`f��c��v�rR�������T��I֪ʌ���������:P�N̜�r�N�E�� p!	���X����_ U�~$�}7����֚ۉ+�w�>l$O�;KG$���le$p\���а)���K�O�x
o�t#mF�FwR�~�D�{@���.��c�>�]�}��fk���p�\>�m����AX��ex��٥�
ƺ{�:��1��`�hw{:�mQ���
4�0m`nB�[�?�9�	��ڃ����� #��Bc�х��o�ǋr��T���:����g����{Zch���:�!�c���(v}� ���О�����S�}p��2���������ͪ�!Bog���	����Oё-4n|�i���9�R��:��5�i�R�]��
FkO!������7N���z8�f�r��'�l�F^n�T֨&���ɴ��-��ՏT�7��&��P0��$�me��~������-��PE5���� F�f�"--7�X"4�������_��X�A���&;�?B;!��~�� ����W�ޯ���!t��=А0m�u��S�N]�@0$�Eo�b��G'<Sx>����V��g kD9�\WH2���ETw6(��;�*/��������fр-qտ�����5[ϲ��دi_���%«��}�1�'t\��L��3<����Wl��-���O*�����M��w�5��-��͑��0b~7�]|I�g��:q�my�ֈ_!�N��3��֔���5�r-��X�.�MLyqA��]��2m��[=�F�|�ՙ�(�� 0��3�)��^�.���W��qw_�H�Y�v�%����@]xY2��kl-�ܓO)��TM&���L@W��;�/������h��'�d���fp&N����@���� X� �
bMr�B�cV���%Z�K�����@ Pt�7�3ĳV�S��d�w�Щ��i�v��M�F���|���3u �>�W3Ga6�D�ZB������sy5YӥQ���͐�ոqGVU��'�/�	 ->{����3���4)�Lt��\��h���`����Q��E^�3"��0��${�B��o_C�"Y�G��?���Ŷ��ލdSD�yŖ�gxY�a�i���>}�@���ᚎ�-rUn+���/V�<䐞bW-��a��A�\�D�6����Q �^���	��8,u�NA��Q��LT[�J@���j��"���V�D	��2:����ݩ9/���[��͑l��/x�Z�?�P��c�E��4��cJ�����?��AF"ڣ-c�Z&5Q�XsJ�C��"v%g `����P�� ��fͰg�f�J"���M0Fh�;����(�&�Y��N�B���|X���h��N;1W�r7(��j�)��>�<l%�y�'Q���'<�-~h�l'wM+���� F��ҥ����T�������"�dR��*[�_-��s���dH�RŦP=]���[#$qvX<:� Oj1�d�j�f~���J�nO�������RcPS�X�k@���?���U�af�C�<��5"�j �Ӈ����;;����q1gL���c��G�{cdcs���1��u���nj�]����:]���3��b�X�8�5y�G���h�ӿ5� X^�DG#^�p�����g�u_�݌�l��������^��t�=e͋��	��ܼ��̄s�-�o*-|Jʙ��<���~j9ǳ[�G�;�q)��}�g&�����T0�V�i8��r�J�LT	 �V�z�����$iP�x��;�jU�y�m����D��z)�����\��P#��1C6k�j37y���_0��=����S�<������X�A��>�O�u�z��HkD6	θ_���|��s���o��c��w�`C�?�%�\�|s�ߑ�Tהղ0��X!a�<T�z�� Z��a	6[�-��o��~���5S�t�֩�KB%�e+q2�9�8eP��eZ̞�QW�<xT %r����\����^~{>~*4�U]4ZǨ�HwPJ9�8������#1��<4bOZ��Ђ�0�Gb�g���%}�;���&�_�{Y�0&�����#_�����ni�����0�JjD����Y�%BL�ʢ6�����w�N}�ڸ�Ŝ�:#��w���H����k�������#�h%M�bj��2t��.�7?�yev`GS���ܘƴ~�\�p��ĚQ�|/��`���[�՟���uO-�;V�+΁��zٚTh����KL ���)ȵ� "����p��~I-yYN1��<��g��#�B�=AT�R�Pc%��snնr||PW�>��P����c�����l��K�O>�Ͷ\���+��nM��	�iKoHRzW�c�bBj��Q���L��.ޘ[�����?��p���[^��	<y=ge�X��r�_�Vf4sY�u���eO�'r"ӫƳ��kG�dB|f�ߦ�c���R3/� {�1X\�i�bU�����!�v�Zx���	j6ϼV�����$��	���r*im��bH>��v<��	⺭a
�Nq���2�%��k�.��:�yv��x�ܐ|����G���}K�7�5N��vO��1"Ɔ�a��$���eip�gC��u����|�O,x骭���!m�2��