XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��2p�	����o�C�����NJ���,����)����w�^m��� }h��>�c�~��S:eL���+r��� �edR��8�j^9߬�ّgw�L��^��GP�ˉ��� �M�ъ��P�T���t�?���-||��z� &b]*-+:k��QuHx���v����H�d@v�nXQy�	�`>�'�B_��|�Ҙ����ab��U!�7�y����QP��Ȱ�Z��⣈��E}J���$	�~���3g�(Cϱ2�>�}VN�̨_�5e�t��P�1�ywA�Me�����n���"�&?$�蟚:���k?Ȍ�E|e�)���	���7?�T���b	b�S�[��t�O�!8��t�0Q���@y2t�~��S6��^�3�(ó�Rp$��z�2鼂�7����]L2`���*=��B������X�����F�ɛ��`B VQ��!��Y����6�ɵe���Z	��L�{g��O�M��ըZ*���7dpZ��P!����t��P����VwRU(� D۽��6i�@l���=�Ɓ1���y�Te������J���z.ύH�(�S_f�X��ܫ��M��_(��!:*5!�"������qq�����9����/A9�<H�ɆgR�I�.|/H��!}Z�ւƴ�=_5��A��/��6�))�F��W�nh-�i鸑��m�Lw�ȏ���1���p�{E�ހ��I�r��>�!�e>�ˎS����Ŀnc�a�/[�8���-����@/1XlxVHYEB    67cc    1570cw
��u|���d�zD/;���7��^�|�w߾�H�����7@� �~�3���Eq�"��2�,���x����PqNj�`
�ʧ���l����Z�l'պ�@D���Ż�^	�}r�N���4�:�˷�h�2��{�;8�tFr�ڊ,30g�'�)��Y�b:|�JyҴ&^stY
�͜fqq�o5��ߧ5�/N���5��|.�����BU�n2��@8wj�9Z��k��+7��wf핤�޴�sQ���Qf��w.<Y?�i)00��>S����׬�wv<�]�v��]f6�Q:�_���­iS@�nb���v�0�lPs�<0 6ݟ$L���$����$���Lc]�n�I��-��5�ɋO�R\���Ӈ�"�C�.���dx�|�M��O^���ILje���bo��v�AhTRz���y��㯟;�z<����[@%�Q�n�<~��!I5y\�K�ch8�",���+��o�#�(�f��j����+�:�%7@���M�0��At߭Q��%g+������Z�����H�t��A���M�PW]�'���7P�o"xƘ����@��k���<�C 	~�K��k͢S.�X-P����%�|#G�z�c�Id��*� +v,J�q���j�v�o�z�Em5��0)<��uj/��N�c
�|���Y� ���1�[�q�7�����a������3���>Z������f�S�2D+2�'�/��S`!kZ���V��x1]?���6�\x��]�Fd�Qd!E��Zy]��ť���7����,}Ǹ��X��Q��{���+L��p��5%����d�67wW�����Tk����ٚ�V���mrV�h�֑�I����"B��25��ݦ3T�WE&����)�M��H� �
<DX	AR-�(i0}Z��Bj�BP+Qi	�D4J��j�S��|AG7�����S��xp�.��a��6�U�.���-_�,}nΡ�B���J���Y���|h>yc�P��4Q���'�H{uy�R&=r�op� 8܀��� � �7E�n�WG2h2��:1w"��1��#���V���a�Q\f�'��S�b��q�{Zs�]Q�l��k�̴��*�m8��f'����3f��*� וi�� %����d`alܬ(�ޯ��5B��]π&��G|^<3�"�]��oש�,��TืEB�>�5bs1R���3��M��0��/��&ؽ�]ojU�v(dl��u1�a���X*�c���y��(�������~��2�逊�ߊ��[�
'-k���E��Q@���^����+^� ��m.��:���cs1���}���F��xC��Q¶��,�8)w�(���?���!�+`��h o0��G�4�hW�-D
�+�k��?�����N�q�.̩\��Vq0.�?���涭�E�(��u���������y�!��`�gOʅ�!E��_F͍�HC�a��ުt��m������?�KP���>���Ijl8��iy4 �M�ϱ�C��^Æ�WU�>>߉��V�/&��Q��RnͱM�X�-Ĳ�)�\��M�;#�凴�P�j�0�����ل�� J]���o�dl_�^��}Yc?`��i���������'��g�~�h�� Ic���Q�ؒ��׼��kTs�eR�C,����s����Y��쑔�^bKM:
�.�[#4����1�2 �����������<��e�NV�5$l�c�H��[�I�nrt+M��MQ��*�@�jz	&�!������L��!���ɥ����MtD�V��կص%�B0���:�z� �=oKP��m����*�OG���|EJX&y�N�P�� {*����}�n�;儬L��͐������J�,��叵���B���zf��]�����w��Ҧ'�#WL�B͖�MDq��"I���ABW��mC��b?��a���>����=�|A�cԪI ���.�[��V'�B����9�Ƙj�;���ro�ξ�by���J�5/�鏄�IUM"�W#?�� 5Eh�8H����r����@�a����# �Z��Q����}�����$���5��FKb�Ѓw��B0���؆d�w�^���\B���[��� ���W�\�,�y�NV��v��a�ri�Z�=��<nf�'H�U~��0�q�r��!��Z�+!*� �'�s���*��/t��(�>�55����\�[Q'��< a�������0�o�~�mGL��E��-�p�9Y���[d��������
.ެ}�v(����_f� w�i�� �#X���h���1�<�������A�;g*�i�ST����P0�7п!�?�S3!���2�f�>Q�S�*A��<-���#2������J����e8o�}E/��?R�xԔ)ڽ=��E��N@�gEZn�mY�R�r��@�
onETw3w��i��i���ݭ�!]g���I'C�?X��?�Lj]�IPx
�W�=�"ѓ�^O�W�(r�����Q�(���W����@Z�b8�;���6 %�Lb�9	4	S-�22Y�]��1��ұlZ�w��)]���L!��-@_�m��R<t�.x� >!)����X>I�8F�v���p��iy�P	}�L~l�L��h>d�z �}�J��^���zn.�5-#�1p��nt�yX��2w?d�����E������Sy���X:�O
~��C~
TS�׭��Ƀg	4�V��W��kP����u�:���ؘ�˒r�gށ9h�
q#�XyQv:L�N��*.�9z�A�a��;;��b�e���j.�N��RZ��Ɂ[���%r�T�w)<B\��������s�j�4���݀�Ms��Q�۩�q��tG���d��F��B!-`���s��KRL�V�rYD��kY��E(�� ��.��09i��<���[���x��"d9p���p��<k5��n�D��>B٧L�O�-�6ɼ����C����]�!�C'����g��0'C��c?����G Z�'f2�99�,�=]�B>�>Z�\�l�����6үl��ѡ%zJ_�U"&r�{���v��.z�)�O)ߌ8�r��\^�P���@����J �D�[۾��{���sÜxW1�8��bVp��b�d_D�^P�;��_�S���&��N�:.�%�
ua9Z�tMZ+�(�z�/���u����p�o�Q2:��mDvN��{���t���f-��;MS伿�Q���l[�`�ۤ~I1�1h��*;.y�9��jX���r������4��+O�:�Ϭ�GS���.&�VY-�\�x�z IbP�ۦ����{��e͉k�D5��}�"���=�@y��x�
͘O�������|Gn��Ϫ���V/�-�H��p�V2�ӊ}�D��>�hn�} 1��62#���oQ�!Ja��q��r+'���Բ��*q��D�4{��߼e�E�d�3� 7�� �6o��Ei���`������k=����A�HZ�b��P�P��׻�^
Q?�N:�xv���:&���}�:�z6.�mڳb{�YxД'�)��w+�!�̊y�Dj�H���&�̻Ff��J�0�wἮx0c'�2dM�+�]�;gR�V�Vi�{���k�Vׂ)�������J��m�x����g����NX8�g���aM:��m[���� ���I���4P�mr��-:�s�[S���٨���������9^L���< �0��30a!�z��ZJ�DN@%����e�5%����O�jhzy�JG�����m�#���Scim����.��s�ξ���{F�0f�?$z�i�%�32!\�%���{��B$�|�r�]M&�� �~*�=������Xnt3��I�@^cl�Z-�XB8������a�)Bz)�\�L
N3�N6/'�5�1s���WC&�[Q����?��,�Xn�xd(-��BL1!��JB�l{�@�&?�zuƪ]�l_?1�����
��l�ƦXKK�i��9��~�C�/M�+Ñ���9d��vg�ȩ=�7UP�ۙ��{f-?�5����2��dThŽx���Ny�}��|R4r��%!�Yw�a!��8��e���?-���~�D���MQ14�R�UڋX���B&x����bZ^sa�1�(U3����B�X����ER��Ү?�f��ݦ���W$2�ٓ��q��k�ج���A����9G����q�O�VN
	��|���"��/^-X�b���3��c:�7��_.�'s��Zo���N���0jk��|�%x������rD~��P����:\ڰ�O�xm��Ys!�����=�b৯N6��Z�M��]���N�U��ޟ	H�zM�"�mŤl3�.�N�/��2�ՖU-��`��X��8y�{��Kt��)��0�[YKN��j\������;���bs=�~�P��o��vm�q�Ћ
xJ�RHT�\���A)Ǻ�(:�_��~�a;k������f.��/Tߪ�&p�:)�窑b�.iy��	�G���"���p�䑠�X�w��C-�3"�z�@�y�b*�I�ص�:��}��>2�n�5b��b֐��c��0!��Q�}�p�vD�r�� 5$���MK���ʻH��{��ѵS�]T��5���ð ��w鞯�o"��G��΍.�VcG�,?S|l����蒲�5�o�ŉ�M��s�Մ��v}�_��/$/f�h��o�����6���Hт����G��ԭ�U���\.�l�1}��rk%�G־&��01��%�E����L�k۶v�-���&J@S\�B$:JCs�ʧ)�_&ڏ���M2AnY�w�[θ1�~�?ƈ}Ph�t!4A퇚��RNk�+̖o\=�r� ����E!����Ɲd�tKeZ����|���tdх��$˩4�݂T��L�LS�jsO������^�f�z����q�*�*~O
+Aդ�On���G��#���w�D|эJ��sW@�!kk�)8���u���J@J�^e��&�g�2��ŀ8`MA�h���� �6'z�T]����$17���8`A^�&9�꿨*�q�Z"�ڎ�}8z����i�B��Ѯ��PK� w���{�	��@��k[�vk=�%x/�}/<��zFlВ���N3Ok�2�O�2����-���j`�km�I�-C�[C9W�a����}uт*z>���%9��i÷�}��#ŋ� \�R3�Mf����Qe@uÉ��d]}4��U2E�~� �����h�y�ߍV�ex��F����kG��= $����M)�βM@Pv���J@3%p	/����u^�9����}ɴQ�`���.����(�
��cw�z~L� 6�>�溗:���D�,�p�a�p(�Ȟ��`��Ά�q(^U�