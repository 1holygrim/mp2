XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����C�/WS<�M��ߖ6�'��I��a��]����gbnF�&�g�w�(T!6`�\G��v)�DS�L�}h����;��?ƈ����-�Nς��(��z����P�%��,�m+�ԥ�l�\`ba�H�tr��w�]��9�œ��lFӵ`��_&`��aO���k7_��.nG �
1��l��w�a����G�$���/�7��kS�π�Y�oG��ϟ��[�H��"W� �o�TI
50�����ܫ��J�ze�K�ǒhQ|�Lm/-gөjK����7��\��r�"��@L�HM��f�Cr^9��q3"���Vx֞�A&<re�0�jf����eM/�Z\`XJ�'�%���%ͯ@w�b�=cS��&$�t ܀~�zW�<�MMJZӗ���B��+�)L�C�-������Q۶�%�%	�2a;0�t#�:=P	=Zt/:�#�Yr'�JRXq�E�xm���PT:���>���&��0mɽnǿt*T$L�/SC�^���۩4��w(��̙���h����H��i��ja�+��I���2�跤w2���2���}n�^o�`)"�q�+�}�R�쿊N>IS����\�2��`4��Co���S�V��(�s0r�8�_�!6�T6���������0h�.���"�Hv�ʳ�@t[�C�@�ɰ`+���6��������݂[������������t$%wj�#�]Mܡ=����Nk))'����T�Q>-x�EL�Y(�;T�s��t�����J~�qXlxVHYEB    fa00    2040nODC�kr~'��`Ť@�RF;���VI�~lhF@1���`�l��i�8E�9���\	��Z{��ZP���@�G{�)�؎Ew��^��Ё7�V3���e�b���U�֭��zus�c4�ܧ5<k�5C5[����j���o;����ԅ5�DoDFdi֛��Ϻ�Me|�o)��sn�Y�J��=T'	�����j��kK7�o�蹰I��t����
�/�r��X@��%l1��7Ӡ%�c�6:#f��s��F@�)���ျ�X#<�K�6�%[p���"�o��iު�E�,��	�D���X�'@+2r�t�]W�!
K��pa��#s<:�b�U�N���ݢA�g���i��1��Jx��M�h��q���w�"dj1���R�<[��nR��E�T�ܿu_���nP�-')�o����B�!�N�O�MP(��.įm�|�y�7;{g�I:\M�W�a���q���陛Upl��yqr`Հ�������������O��J���v�#K7�N�il�5���d��@$�[Xĭ��r@c��%^Np�*��^u�>�却p�"�8�"�g��?��U-�WH���֏�KO���H�odK4�4O>��N,?$�,�
7��=��������A��4�x�=6��_�Ɋ���7��AV���;ε�4g�Gh�?��6(?-pN�b:)t��G5f��z86T6��)��[I��9���HG�>E���+/����������8D�2Hs�GdKJ%�O���\���&<M�����ȵA���Mŭ趙J���U!�JE�#�6��0ZT�	���h���X`�J�Q=�Uo����6��%{���93W��ΰo��w<�g�9˰�&�lW�DR�N�4(.^���Z,~�-3�iW�n��{||&5� !{���09*^%/PV�
 i���Fn������d1�ۃ̚@CgA�KUP-@��pb��T�½#��DI��aR' R�<�;3�"�qQ˛M3G�%
%�(7�2xk���:�I�7G��:�&�v�ω2+��!0��x�0ޭz�&���cӰŉ�Ѯ��4c��EAn]�9��L�;�h�)p��s���@?;�De~čYZ����L�Y=�fE���]8h_V8� &���E#�����Ut��'�Ѣ�d	�:��� �Uz���u��ab����-1lIJ�7Ң�܇�}O5Ͷ��5�,'?��ɤ�ϖUt���������C�_�Ld(�/tG7�x������#t��0�B u;>��`�o�5��㠿q{'�3 n`�n�Hi����i�}U� 4�����2w�ė"y���9^+{'�w�=>?��so���Ep̼�ٕ�����-�J1"�3�Fë��-���țTQ(����Qp��4*$���`�?3� ®Cc�n_�$�&�\���l�?�8��@L`%XrD��kL��Н&*G�wK���v'�O�k��?N��\}wQ�_�(���C�g��-��y� �4+:n8�mgm���GJ����ɵ۟���T�Gk����s��Z�����Ń��Y�a�2ʅmm�랏|�?���Qnܽ��M��\�����h_r�z %і���;s�I�M6H��8zN�'���Wj�^���^�v�tJi[������Y&��(p��ɽ,�i*�H������C3Ĺ~|7A��q*Hr�榞�tj1��J�)�)�F�Ҭ�q��"���S$mX�1�aNC��l��Xm[g�%���Ρ�����ֺ'Z�y�
�L�o è��w0�@�.�M���<�?�(��.��3��S?�����x�Υzi���Ҥz{�CӠE�3�J��>�N�u/Zuʚ"> 6&( 6���䙼�V�DG�����3��#ƺ�%Jnɂdb=�#⳿�ƍ���4.��X��޺��{՗����,7&��:{o1F$%�{@#�%*0�G4{w!6��!f��j�ϸC߫�r2�lE���,�������R�-�s4zz�M���R���W���N�&yU��R7c�=�Ȼ��[P�m����Z��� ���Ѭ7>u�LPH�M��s��PB|@S�6>5b���M%*�����MG�:B���i�~(I:�?�6���/�e�#7��A�-O�$��j��XQ���ƭ���^=`�U��X�<���򃥏^�\�O D_ɛD�L���c��H��t���:' ����������,�0&�L�Tw-����b�|�/d�]	�H���C����4��Pz������Ҧ�tA�2�0R�"���w�O9�ڹ�&��M�������h<�a��Dt�J = �&bi	0����U"|�5?��~Gb5����K�ba׌���V	e�?oXKW� sVҰ�]��^�����\���a�(�ڨRi��
ƍ�w�����@����p�!�g�������&�2R�Ʒ�e�����j�먣y��|F%�=p �v�
8u��{�_��`n*I�|�[��z�-���Z�'�����r|+ʈ���#��"ܓ��n�f�<E��m�QQ��J�FNpꏻ�3j������k�w|n=n�LH��_��Ë=h�!\`l�u���m{���ȿ�����b(?��5�E��>h)�pMgN�
ܷj�v��'���tz#�:g#��-���|E~��f������F�<bI�Qnv�w kL'��Z�V3�z9�Gۗ<�?�m4GI���FX�3AX��p�44w��,Ʃ"X���!�!��>>"qe�+�L��c4VY�M��.�Vk��H_��pA���u��#� A�b-ؽ�i�S�����G��_  ���2d�Y�P	�/�c�e:�,���{�DM���z���9�_�h�}�e-�4?��ˋ=����"IUw�[W����!Z6X�P@�q�	�k��!��sX��l�ّ���s���"#�K�jB�rЍ�u��������:$8#2۽=w�U
Y�J��dAFH�Xu�NM�<z��W�):�n�;�N4W�#�/I>�ϘX�d<	���Ĩ7Cj���Y(�c[�yÑy �(P�<��0~����D�y(׈Oa���Z�)�O�_�R�9�^�!O�����ܬl���>A<M������1�-�f�3n�q�����x�X�/����;��֕f�\��ǐ'���a
�M�A_�x'�W ��	�-j��,���FS�mG����x,̛� +� ksaa���s�8<���d�F��x���2��)9[k�� w]�����rG���0��V)�2�M�Luܹ2GrB���c������H:cU��G�$Fw�1&R�&�S�\n�d�
��{ڢ"�[��3�P�B��J��R��|��ٲ�S@B�\3�gA,w�H�@.3�2O)Zr.��0�Զ[�9�$���T?��Z`]OK��	�,�L���G�Y�����difV�G	{:�''q�-��Q<9�W��8|�!��CA����� ����y~�Ӊ��ʴ�"R���K6�[D�qe�	-���"
�� }�n�No�a���&xU�S�8`�׾5	.�����5�����4�}�ֽ���Y^��
 �ײ�r���?k��ˤ��� )�t�6�R��~��u�u�:)X�;�z���GZ"�$_^�P�A�%Ka����{���"��-J���E�m��WMb��&�[�l���C���*`�}�(�A�(G����Z3T�!�}�;�k�D�g��9&�.��Fݬ	1��[�	�wݴ�~T���ԇ��.����~�]��u��wI�^a�f�b|t�ÿ]��E[8rݣ�zF��B<C����a�p,7΍މ�6��$�)ZVl^����SnIV��؍^^�j����~�+�ŀ`���hv����ר���7Ǡ�:�3�� �jpqzQ���'_wI�;e��.8tP��3�h<�=�S���������2��
�Q@tFf��/$=1�%f�� �t��/�BτVk�@�ߓň��bJ�z��뤬 Ẃ�`4�I#A���gmĘ21��_"E��5����" �^�<���x-2�M��c��%�%I�j�\������t�rꇕm\a�%Z���Z{��޳E�P��I��B&�#N=��{N�N�գ��c�`� �?͋`mIb�v��Z�lb)cK��a$�_n�	:tOX⇍j2΃b�Ж�<��9�>>�t�xf�"�Fƾ���/n5v�Wn��VF��0\�֊�/Ϟ�S��:���%�����0�n�N_���������l���<���'���,��Cp+�U���\5�`/��\h���tɹ��;l���N���u���2LF���4z�fŞC�=O@n3����3�����)�D�����b����W�� ��"�V��q>����A�,n#5kFݯ�ˀˎ/D��C�S³t�֒������Y:����2#�Y�*Ü�[vk��
kfZf�[;Y�ȗ���S�]ٿ�s闲4-�յu .�1~,��b���(g���n��7��i��C���Ɖ��` �H5��d����c�N�ֽS�}"(�~�!���+�雿QelG��ޗ$]�DJ�����WZ�·I|d�wķ��:��HBHY��-�+>�V����S{���Z�l�i��P�N�{AS/~�,qa��jQ3�1���#�A���T7*�WD�"�4�-O ��`޼�룕��t~�ɴƖ#�ތ�6�gpr�}4�!��oxnj�C�ս�vO!�kQ	�d,�10/+�}������Bp:qo��L�ɓ����F�ܒӧMZP����Z��j
�����f���T�С-��Ƹ�&��Q�|�+̳i�Zڀ.[�9w(U�z�Ȃ\L@�a(I��H�.zK,NN�g������`�HK1(�/M9��&���Cܷ)��kݛf��0�m]�o���n(sG���|Q��7�8�hd�F�D:gZ�;��>Z���Iۆo����I��4�MK��>�	t�	����N�h�*�&M��i��`?��Sܑ�_���@������+�ΩUNg���(�O���3�Z���+�d�ͯәSձK��+�0e s��L^��H,�����\��p;��{�eT*����G�݈���D�kyi~�&����L)�C�_b;HHb��E'N�|������>�9�ޔl��ۈ]����ؽ�J7n�7���f�9%���n��;��X6h�Ż&	�Y~�}�xZ�����G�L;X�T�R L�Bbda �VNZ���1�![�-]��I�Wl�q6S���d�_�UXB��ה0"x-n�˅w�U�:z'���!���FO���Ұjs,%��Ky��-�ҏQ�F�@r�̹�h�h,�"������b�Zߋ�h]A<=��G�~�5� 7j��i�$��v9LaPޣ�����wfu1'-��f%|1�?$?���e>[��<������so�]�.>����O�<?�AG�����|m�5���E~���>�c��:�� ��P?Mf`Υ�Qp�T;�c �[�����	�Q�7Z��x	��6o�b��Y�t�$i�U���@����O���5$������5 ���&����_X�l�p��)������N<���zB Ҟ������CRW2���XH���7��ZX��=��e�͛�oQ�>j1�m�TS�~�o��q/��F3`���.�����嚴Gi"bޫ�ݶ�EZh�9�;q�"��$��Z,���lc�����'��aB��5
�y�榕a$�笺�qU;�����=���O������j|.p���'0*J��٭z��=U"Z4������p{xHт:����^^�-�Y��'fY4�7`�@�T��N�"�k~O6�m_[e;e��rBFt����¤�N���[z]o�23Z�v�D</�!A׾fe~���q�,�IO��%
�1{������kc��)�J�����/|J��FT�T��<ǟqY]�$	n�ݨ{�c�=5��&�s 6G\6m�����F���7$~��h�C�O��)��h�,6m���Z��y� 5y�)�Y=�oķ����ݍ>+LĢ�d<NQ�\B��Q��6��7c�iL�܇���o[���x�>�_�sW���D�ǣ1/�٦)��t�!�������{B�H����Q@��ð��C�K�m���%1�8�l�!���'&��Q�Cz?�N��y�%�|�jz�mdP�hx�ע5�ldM8�wO�vH�����'��n�[G��LN����q� ɤ�K�º��!��C&6�"��az���"+�����Ol7w���B�H�m����5s
e�m�ũFA��3�~[dQ���\��T)�x�|������|�
8S=`RSj��&� ��	�o�	j2�F.�Å�.��D�^Z �ފ���|�.�sG��D#�l���39�x��
,���b�q��87[�&|����� ���Tň�qCC���sCNd� b5U�`�(i^�837֣I�V�I!l� �Ɛ���&޿Dw�2���s�??�dZ}�7A?����SцY��L�}������y���*?����vA�N�e (ﴊY(F�<�L�vJ٥����A����nd��-�Z���
�����c3`���n���M�K�X�W���#cDq��R`�A�V��w��WA{�����yb�-�;4��#��mG���(PZ�~���i7��8l4dt<�sS�˩���.�A)�ƞξ]*q`��< �#o�p��rbܼ}�[��Z��W/`j2���S���ؿ37�LK=�M4p�`-�/4�+wZ8��zǤG^��7��6����X�ʓ[�9�>C�9����r����3�}Op~3핗�u�)���?����o���S�������[�{�����S#�y���S��D�ˊ�(�����*�`���-�!�`��NH����u򟃹Ō�A���s�-N4�Cة�N�+N�wc�+���Aw�ct[CI���@����A�4V$�i����Ԟjnt���,Ac��Ǵ�P�[)v6�&k�i~D{�ξ�)�Ni�7^�(�s����Y@9\݄�:����.�ۨ�d>��ץל�L�`�b�̾
G$��	m��(��h~%�5^�/����ǋ?��l��-��{�nx*ru�u�:�C�l�YlT>��	����]�ea��PQ�+��=�h�o���𘊅�}�h�f>Y7�E�@�ߋ��Į�SL���T�0P�;�s�*�D��M�\�2��(�)o=�\����Y�\��E�奺2��&�摸��r��! `����T�L���3�_����2������Clώ��g�OYQ>F����K��PD1Δ�|L�DϹ��7e0}���jj�A�������km
���±n�ϊ��*��#��4��U�Bz�nY��F�u_f�E�d�-��;x���9Rm�f�7|s; �UA5}L�p��sH�����w$2 �+&ӳ��V�L�JI���uy��Q��P��&�07���L���%����5�Î!K�r�e��E��t���zpWD��f��4�B"E���vxB�G4!qG艂�&eTC� m6�'��(F!���؈�_Τ���Χ"hT�X��)GU>��I-�Fμp���\��`��r5��> �I���P}�	H����F�'�is��
ڷ_�|a�0�~��
��N�_��h*�;�P�s�,�uփ����[�`�K�8<aWb��I��龏vM�j{��[�iiԏ�����1��O������p6H*�^O������<e��/�@��Kcc�T��KMo+��qMt�PQ#}-|h��Qo=�6�pLO�*�4����$d�����6k#��cG�[���'��m�� �)7��X��W6b���tn�-c���;�ө4$ΜV8�#¢�-:`}����/B5p�v��{i="x��I���#��ǮU}J��0�����T&EV3�$I�wayŷ��tIk��:�VeyّGJn��q�gϥ�V�v�u�g�-��{����ʌ�LU���A}�	�dn�*��y�:�S�pc#kAER�ƭ5��R�\�������u�XQX��&��7��	)0)x5`�7h��QF?�XlxVHYEB    4f62     b50�u��������"��4 �
N�O��\2F{DN�_}xe�˰3�ŇaW�|���'c�r-eۜ@���<��J�o5C��N�Ղk9T<:��B�+ӺJ�ͦ�$�E {��f�+���%+"��K����ߤ��v�����#�r{�(�x���H�o���O�{P����d����:uX�	<U�H|0>S����^Y S@1��UtUp(�6��l��R�4=-a�r�8���{=edO�$�J��+��H	��I���ʆ��Mn��`�����ė�6��u�x]�&�F��$��ie��
���i�Mf�=�}:c��CD5<�o�T��B!U�~��w�P�I��׹1�g|�ᴅ�}+j�#�5��Z���ЂZI�$L��!��t����IbO��pM 5eS��$�D;4�����i"���9
k�J(B��0�S!"�d�
��'+AwUԘ;�0�Um@�,��Nd� �s�Z ���z��#^�\n���	����!�p �C��N0�a�A!#��Sc��5SW��eH2� �\4�Ol����� ��B�KVfL1��3Ł\�"?wg!�0�$_��T�֊!���P�}TYn�g/G؛!F_��
��×���B��P�M7��$�_؜�|�R`�f�Ƈ3�3�aH�t����������ÕP�	2���f/���Ys����kyυ��~8��j>�2O٢w��ql�rD�_.j/�)>#	k0��O�Ժ� ��V�wj�,�bj\a~�����~�P0�r���~�4b�{J��y���@�7�r��G�"�I6��C~�C�r{qb���r8͵�OCS�4�ձ6��ĕ���R2Rm��C������g��:W3jyL��u]�}�h�Y
~ǅ�ʰ�|^#�k6D���س�	�����p{S��M-!�ڧ#]��L1&<��4���� _	��|S��[G�zFk�0���`ԮC��}F6��-��V�Gb=/�UD��ł�U#��+�}��;��ً�-F60.���z��h_����9s}C���!��C^�9qF�	n��I ��[虆k���q)�)�� c�%E�@���'?��3�h���xs����{s�5��).�N`A:O�d��X㗰���vȦpą�8E-�%A�EZ�3t뜏��琱J��::��������</��KP�<=�`>đ�אł7�h����IۆS"l͸py�Π䮎w���r�Ϊ�|ɹ=���k_�{C{wH�Mïeu̲���S�� �3]�� _�ۆY����,q��(�/ل����\�~��-�q-(�l!�Xo<;W"���T���x������{(�-��U�� �h#7�6�7J��B�Iրʮ�J�JW�f�h���Atҳ� ��@x$)��AɈ���f8�G�R�� ��VFeX.[��G�ʁ�~�ϒa��"Q&�l3I �O���A���?]=N�x�!A��k�<���J���-��sU�e���6�0�_�aL(E$�w�Q�&h=���clA�x��\v�����f�w��w��5����A�86������ey7M��`�I����&��L@O�U;W���Mn�vn�]2Cj��s6X�d�Q�0��!����0�p%��ax�Ό�NP�e)�c��j��b缆�[����r��G�w�5��@���W��;�ꥬZwt�&��O$�o�,�qxd_N^�:K���Y��"VM��b�)�#�Ns�Sé!u�����ok�"v�����+ �K'�(�I8��%~����FAM�)�x���J�%�='}����Kl�ؾ�?~�pi��0�Fγ�aC��D�A*��-��YT5-n�G>O��:#� ���~���_j��C�Y&��#���h������3�q�0�F$	�ZH�hu��%�V�=E�] ��͋c�T�X���:��ѩ��I���B^���2"����Sݩ����m������1��g˂�v.���0�K'��|api�E���֫Q��?�� VA��O�4��=� \x(r<�m'�WE����4]t3|�w��fh��4�3�"�n����ES�޷�!�T�qQG
M��C�
}�6s�bQT�GG���d�3�;ao�t�u���0M4�m-2~��Bz6�iR���s#Lyg�x��)��t'�Eb��7�_�o��Ǽ,��!*b^$�LYh�#�[��>4y�������h����@��:�(ϳO�2��/`O�}���T���pΒFN���p�Ȍ*L�@*���ʟ\f������[u`䋪�?�m��ĕ���C��o�*%=G,��m3�֨1j�2`�B����$�PRj�P��~�]/da�F��1*��!�����<<�6V����`E����?5!��:�Bk6�S�xh�ڕ`p+v�+XT�<|��En�z�����W����9��a���t��]�l�n�W	�Yi%���9	w�1''���Bm�^+�N\"Ս᷶^y��� �
Oz)<}��M�xG�~X	9%q�P�3�ia�7uL�>�GV:��"�[��-N��}$�p"b�1�k��^S��ݥ����3���i���<SK��܅�^��ȑ�Ύ��� c]���ʭ�¥\6@��s��r|H�-�E� \��Zi���-,��nL���p�@��d�(H�E��l���F}�V����Ѓ�oPo�Q,[�J���ƇAi���`�l{�m�� Bq��%�ټ6�0�+r6`)��r�A���;�)G���Σ�eN�eye�('�P��	��ko��5�'�`N �S�-��n�<U_���!_)9��I.�?�$���՘��c���