XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����5��6�h�GSS�!@膴�t~�)A��	U�խ��2A$��\�Y�_��[wu��������_�nG�<�e����!��v%�mD G��NTMk�QͰiѳ�!�&�ᡭ��"s�N����;�(��q䃏-8�k�q^��m���KEP����,�b�
:��|�C�`N�4݌@a�Z���'�����8���U��6�C�xsD����$��	��]0��9]G��6I�;��"��&��Ǒ�姥���G�I��>�8�;���c ɡp���F<CQ�8'ι�dӍO+7�V��	�K��"�t�뛽e+���=���7Q�x��N!��Ei�x` �G6|�g_��˼?<���o��]��:F�$Ȓ�� ��4<4�d���A�������Ik��^E�� 4^�Z�[�5����_��p�\�e���u1��,Esh�-8�ޒG�0bJ��Z�.��޾�?Bݕ8v��3�y�ue��CZ��|�hE �-�\ׅ��@7�f��L�6������\.}})$h��G�ۛ���x E�^z�za��SJAT��%�O�zmm�ٸ���H����@�]fѢO9|0�j�ﭓE��OE�y�5�E�8�tITÛv^�z]�+b�e~�o��@B�:	9222?�:b�n�?S��_a���c9a�U�>�T��y���F=x?g�����쪪�S��m����4>�a>8`Y���ŉ1���K��J2wJ��hչYl���R14�x��5�wqS�N��U�F�XlxVHYEB    266e     ad0�5���7>��~�����RF��5]�q�x�s��,�Ԑ
'^n��g6f����7��.$c�/�h"]���� cye3y��aե��Eɤ X7�����}C�s���lt&R��jv��u��(�x7%`^�!p�ǽ6�FOD�g!S�n��\a(&����.���ܿ���5�t>����:0�
�P��JD�Ɂ��L�~qk��p����>zK�n$������&2<�2�W2����W+�Ln��_[?�� ��v�<�WsA������Q.
�m�a%�֖d�a�V�'#��yE0��ߌi��&'o���k	�=�>�����_�:�f,��PV����&(V��a�P�E���{�<�O�Ο�_���`�g�N���-gҨ�����y��\ Ȇ�o�bn�L�z�'��ڷ�$3$�s�U��mc�x[�D�[)�� \w��q"OZv��}��BD�,(�g�_�Z��U`��&c�t�����An����@RO��H7�x�~���/p:=Ә���e)����f<����QHΖ3�M!�rR�>A�"�1��)����A�3�d�"�$�s$ɦ_� >�IFp����e�����s�CO	]��xS�kC�Z�ۆ08y�9���'+]���W��4�o�J��>P/f�K]�-f�}��Y�c4��ay����T��V�>(��ɱU��y.oX�ud����X�"��V�d[OgK�EF�0$F�AC���V���ǘ�,��* [Gy���3�n*_ɐk�0�����I����V~>j:�q�Nd�4�-H'є�i�-��o�!o�7a������"'��7��8�����j��\n?���wf�L� {��/Ws��{�r;�nI�����r&�G�R��ګe�u��ϊ�����O��P��Ͽ�'���#h�"�(�	�7�	]��jz�.W��@��O�;�<�lp���m�Q�/	�X���z��Zzf�*A9�J���7��ϡ�R3��0��䮸�8�;�v��4�$��%y<��rc�tN��(9�,��oc��\��?��lG��M[�<	�SZs��|+�A�Z��74J�U�i4ś{7����.�_{�A1Hlz�N0=�$I�{|�{7�H1��o�7'��ż���E����OP��P���&�~�]_*JK�(нp4�A��4��e/b]/ ������B���Ԉq��n�X�m��/�r��{���Ԕ�Y��G�a3�(߫��n?��#z}#:.Esݸ�����]��A?��A���vY�?c�Qw\Ķ������܉jkM���<���܃6�Y�8�x��{���ൔCB֨(��A�H�4�1-�n��ĭ`�"��^n�g�Z�Z�Y�գ�������b><��xg8��1��"�x�_-N������8J����"yP�ڶ%��Y��Qb�`]B�!f��0�9ݝ�����'�+�G�k,^-B��b+^,*q�2�<�C���`�4��#���7~n��jmW��s�'I4�W�X ��H���T��������	�E���������X��/�ҡn�8,�n��n}��>FmU��9�X
�������-��O$�y}�L	<�(C��3�\ıK���Q$N������t�e��5�K�^���L-8yͧ��@�?���τ�� ~'2�{�3A��gv�h�E�}Zw���S{@4캙^����v-#;�����ҿA�y���Kh2O�)j���s�/��@����:���YƵ� ��p�>��zN�y=�R%�3H8вs��r`�
XS�Ŀ ��=��>Sؔ�.�� .�ݗ\��o��ҟ&��qp{�p}��=�U�������+,�S������e�(@�8��-�8V*n^���"�ѿ����.�hAh�؄p��= D9~�Kj5�ͪ�Ó,���5���V)D��o�3+�w���;�<�z��,�͑��G|,�X��g�FV��K�����L��;�uc]S:��b#��D�K!+���-_��ko�q�������XG��+����S�P'%�LA��ep}5����t~G��W����d�r�?�u[��@�G���H��qE�� �����c�d�z����lR׏nYmJ%�U2vl��9�fW�dr��������R��fDk��h���:��V�'�I��o����ig��Ѯ�㤈��z���j�EH���6�2W��	�➪\��ߙ}�� {b�����g��LW��<D&��t�W����j�Vwe����lN%���`�$���^�b[��@����ބT���uJ�J
��!��9)駒US�����F��a�}�vzm�Z�G��NE)�=�8m��C�ȧ�[@;�˿�hI͜��$d	WM"}u_gl��� E@[������ER72P�%7^�ۆ�3�F"���[��=-,am�	�6�x5t^�9r�����㎭���[1j�6'�����ކ��g������O��Odק����O���"�S�x�y[�-e�]����"���^g��~�¿�OM�f�$�>� �Oc�,���vfs�q��A��UR!h����V�G��@3'x����}���u�,�Be��F-��-#^h�LD�Z37e`G7�ꪫ}y�"��%͢�=��)���2Ay���j@A�_�$�Hp6���",B��s�áhѢ��Se}�o��8����@�����W���+�^Iɇ�_�H�I1�"��>+�