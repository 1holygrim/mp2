XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����b�٘�9ڪa�V���4�G�NIM���ܨ�;�����^'ܣ���1ٖAJK� x�ggOuڍ�.#Y�����}��M�R�岮���t.w������w��)�FO����cJ��	7
�\=��ě:�M���kS4�|���o�5vŲw�z5M'����x�o��v��*�O����-'Fr���w�@֛&�V�z=�lL��$�z�?���[�����L��-����P�Vt���p<|! '�E�o-\�tYZYe��Se��s���[���
�v �Ć�����y#���Ĝ��k����ը	��Ikt�����wZF�=.����5]"Oi%�����@��q��"Ƅ�Ɉ��JBRvk�^��c�����y"u��,�&Ըc��ab�Y|�W^�����P���q1JT�D�'��ѱQ�0�
rXX�U���e�&X?e�jz�8�E�1J9���Ƌ+P�� ��咕I̊g^}���S3l�g���^]Wप�h�X��<�O"gy� �*r�8E��;�e��ww��Ԡ{6���'D[Thl6b�3
S��	N����Јt,]���6�8��ѹ��{������������0�1����_�P;���	��W�_!駞�O���،�é�2��)A(}��X����Ѣ���W哇�3�J0+'d�Y��(X��=T���DG��g,�P�����r
�z�l���J�@����Q���F��6�	ث6��-u�0�+e>�XlxVHYEB    95d3    18d0�<�a:���\ߍU�c�p�.+���"H0�Y����~����IQ��P㫻��+C�U*���R9�g@����tb��y��?��XN�eQ<<�Q(��8�e�������ץ��!%;�p� �h�Nd�����}�L*7Q�2�3��0�*��� *Ra��b�4d,eg>�EH���H�O�wYw��L�E�C�Kρ���@��fY����\����l�od�s��
9�ޢ<�4�p*H���R,�W�����y-Q�Z�@� /Z��v[p�2��1�tsW�X�5����)H6��Q�=A���r�e�:�P��v�>xӗ���b;���	�ԜJ⪘ҩsY<�h�`�K�P���8I<b1���ι����G�=N�1c�*�E/B"��H3&8]�O^�_���m7�U�n�����u�ۂ�)����E�Ȣ#O*��y�[�ܴ��_�CV�M��z-�f�xd�n7UY�0�#����G��ol��W>���͉΁~K��r~�l���6�����ǯrɞg�H(����8Ƕ8{D�[��'@A��^��?_�u!s����ggI}4|����︦]b_ ٵ��91�N�EO�"��oɩ��7�.�&|9d��QΦ- �[��|�Z���T0��q�������61��x��<\�B��uZS��#D
���:u�r��ߨi���8_2����ڼ �a@is@�k��3Fų�DG4��P���vʖ�?� =ĞOы�>l���c�\�Ċ��A1��Ƈ]�ay&�>�? �{&��;�Q�(g�uV�ﲙyZ ���m��
H�!���yx��]�>��W�1�a�#��P��y����ю�b$0U���I0�������Q6�](s�N�{�?�3r�F"T��(;R��!i�ggӢ��jA0�}��_9��Mӄ{����]?�8�`�$��	�O��P*rhf�"�%͡��+�`y�5.vٝ&���w�*O霸�TF���Ÿ/������|����O+�R�h`�޹�wYk+���v���G�P n��G�=�D u��9~R��<�tb
����=�o>\7��͝^��d+V� �s��?�'�@|w7�1]�� �b�
$Gs�q��( �)t &R*�Usf9N��(��r�R�$��^+��|z���) K=ia�DK2�FQ�E�ūPw�F`*��u��._0jz�_#�%������]��_.�u%g�qO�2 D.�ˈ�̾�#���tu�I�S�2�� ��@�'�}5^HA�")�n�r34���i���$���p��J��SM��]�N�l�1�zB�?r��%L�ɿbe��x��8Vs�f��Ly[H �ӽ�|�n��g5Ƅj�Zb*"�+^|��|'ţ�>��rg�<)9�6�]�K̷QL��$��S�PO��8r��s5>�:�'�ؿ�����I
��4p8XFx��J�?�}�C��*�0�t�?*����C]�g�HC�.l*bO:��E�Qx�+�Gݠ��H�Hm�����yj/�w�M���Q>~�'�h�3��z�͕&��61q�H�7���i�*�p���,��[���s�.ٙ�ԯ^
�.�`�[�vҺ{�e;�)�1,�]Z�:� �쓼���7��Pe=��^��\^��W���I00P���_���>�A�n�xt���u}3L�0��G�X�p�����DX�2�6��;�ϡ���L��ލ/�3ޡؕV�޺0r�rsj}�d-��Q�-+t���l�_(�]Q�6���������@|�j[�9�\epy�����	C�=���%���*ެ]A�j?C�M:cu�e0I�<�J^��`E��xF�y��I>�p J67��jI�j	c.���HX��������G���^���!�K�m+C��ګ����"�)T�z��I��$��U�%��:7��fH"�Y�bHN���r`��&I:[�}-\B[�D#��UĠǡ)���j+�{�R��v֝�D��)ng��h��s�\�����c�af�+�i�����e����aԆ9VׯUE%҇��>�r,��3q����mV��=�Ҿ��p\f1�ff|}��<(E�?� �o�o҇��L�Y%���>���|��w�,S��~�6��;re�JXbyp�����9yї��/Rbx��c��S💟7�[���[=n��´R��S���jS�.Oӈ�ru9��"�=�i�����dfM��ɱ�k�,��n����wሕY֤M�-2x��+���� ��`�T�Z���ɤ��~��s�iZ;	�h�_2ÑMQ'|���<]g���W)�<EʨZ��
�K��M���ʴ0�y���k����������9�XցFIA�[~�H��0���qB�z`m��A���Sɣ�@i�"p�����s��H�:M��{�gj��Ɵ��F �6]D�3Ћ� ,.�&�(<&�bt��,��|����{_=eZ����ف��������	���\�%?bN5�^rL��*�e#g"��'��ݥƤ#���<(��C�+�"u�ĔK�G3{Apn_�D��)T(�] Cq���]��ۭ� �^V�R�S��(�Q�th�8*���
/���#���J��|�k�D`_D�O��j�u3��0�:��o�����+O"��p#����b}@vB�^u7���ǝ�qeچ���Q�������B�u�0�o��(�T�27=o�|�����gn}?g4��'���ar:�	�/b���	?[~�LW���u�p��j$�\]���l6�q�,j,�c(h4��4�dy��e}�o�}���
�T/)6B9�߂m�`"8�!c��j�)�|�m��-*��&��FQ_���ўF}q�*e�ѹ'�������v[kosr��r����9�-�_P��֨��S�e���C�7���Ӡ�?h��!��h��B�9�%J����1eA{���H�����۟p`�O9���zM~`G��6L�n�ŒFA��W<r���_&������<sF�UE	x{��r<f;�aK�j{�e	���� ��s���\Jj�߬���FUN �ȍiU ���n�0�E�Ҁ�>�ef�q����EAO��o6�mK �Y�+�;bRL�X\B~��(@=�@qڢ�}O�&ݲnFݻWG�s���`�Ո������I�z}�y��-�+_�I~��,��Lp���ˁg��"Y/�i4[g|^#�E)j�pX��7��S17b�6e���q%��wM*�%�xg)R��'������և�J� �:�©���NTO�����)��~E�l��̆ݾ�/���?e/"���#L|0}nH�e�D���P����W
"Exϝ�zቘ���*\�,�ĸ޲��?�NQ97�E��x_� ����/}�|ImL/���w�$9.G��͔�1e4S��w`�{�F�IIl]6�.�!�� ��w`k����,��~Q��7r�S�����6�3%$p�;!2�?�G�E�역H4��7�|���i�N�|#ʝ#�@���ʯ+�㟒�GBǗ��Ɵ8�Ų:�1���
�f����C	e�nb����gI�<�_�F�ǯ5*� �ć���kA��HIy(��_����$��Iuه{�`�sj�X��	�
�q���%X��p��H}/�f�N��v�� (yv�e<�a7oo�E��8���_w����cN�z�!|�[xD�z5C`�T-�m<�`����(��~�ۙ�nr(u�5@Ex��hA}�$��-/�-5O�塩_�0B@-��fؓY��Is���+��q�i8�<?@�fS�y1!�e��(��h���*�Sj��l\��`���WUP�<��˭����xk
�y�-��E� �рCby;$E��W�>�o�bl��50�DGd�>X=H���U�ɟ�j�F���i����Rb�/�'"�`�Ӎ!323zN%+KճI,� ��G�z���W�M��SJ�0SeЗe_5֜+�}A��mh��u�
fw�rH�(-�y1S4�q"�j��L^������ӝ�Eܞ�+8��W['ɣ�Ϋ��^/��K�έ��F⟻Wf�ie�T��*��dm�0�/���3��	ҍg�H}4hZ:ގy�Ӊ�Б�/X��ZdҝxA~��M��L��ܼ*�.�O�_��Q�F�8�88�75����ˈ��:	W��R �[䀰��=�nEx��
4�-a���������Zu�"A[l4��Sd�D� ��8
��bY!��U���*����UQ��L$����{� fX73c�bN�H��y琸Ep9�N��D��� ���g6\���i׊�Ar֕��nu7v�ŉMS�.�N�-��I)�F��A�I$בF��xX>��tص�\��J����^���W�}�qEt����@��˙���ʹ/ę#sn�3�U��8����O�hQuΪT��[?m>�.cV���*J�~��҇&�믷��u�N��q�V�5��������l$�+�j�mDtu��=�&��rǼ�/�.�b�v���+�����'�����\ZU}�ҫ���k�>O�!��w�w�}u�Ꮎ����dERN���
!tw��\ܭ�.����1�"0�������*;�B���X�݊��;�gʤ�a�r
��^Z+�I�e����=L������X{o�����U��ܧxʩ&���eb����,\��5��
=���0�C��!Hb�D��V�O��/�W\�R�>n����@ɬ�f֜�1��M�{1_g&�O�)��~�Y&�a:Q�e((���m�D��]7A�z�)�T_��2c�����<ʪnG�!�޹}Ĕ[Nͅ����ߪZy��9�ٍ��Dv{*e�x ���g���x�����~��\H�-���A%��7H�q��[��9�hS7	�ϣ�F-%��mq��m(j,'M��آl��ݛ֎F(y�p���572v�a��oL}8S2�n9��I�N��g�@��P�dFd�@�q�V`1�G���.۝/�z�:I�}%�{��c��/^�靅]�1դcx:'�O��Y�M8�%Q�G��9��5S=���"z~��儡W�����KH{67�[��-O�b��)�x9��q�!b�ǕA}�g��ә��ӿ?��l���-���.:�/U��m���yZ�� ��{�\ďآv�A:Q.���Q�7$y��L����uD��e^�sۦ�^�[7���oW͚k�\/�3~�}�� �X�+��������:~o3fd� T�ߊ\0A�ʮ?I��N᭙�R�� ��dW��{L� 	}k�e�[��V���Ըl'��Mg�����h���������� r�]�&�ȃk�qE�o3�6��E,�V���.d�K؛_�:��Z��JvMf~2E�m�6��J��b$��+Uk�N�tx���!��`G��CѲ:(�AU�j3��}�W��c���짠�H�>�����G� �هB�lx�(l �O�v )mZY���k~�-��z��m-s0M���LM�e���g�9uڷ�d�O��N+�:t�&H�Փ1k��~iUT"1�*�gd�䶞�O&�y�Ŷ���\z���3"���`�d��ۘ�?M��CiH�I�P���Q���2� 9�e��f7-����i,u�8��"Lx�0���H�Q���7K�3(���͍��%�KjW�P�wf:C�qP����'q��+��	ȑ�6�jg˭�X�q`g��c�zؐ12����9�3FD!'�Wp������'w���8^4�]�I��	�c�B�E�:�Mo���ո�C�,�C�^�Gߥ��~�%#�b8�/�1{�l/���T���sk�U,γЗs��g�Q�Y6��<BVS���&@�9�Rq�τo����t�ּ��ƶKʅ{��	��v]��r����T�R�n�������o��_?������HO�3:�؞�9�����r��E�a�T�ve�G��#�eq�Q)�&���Q0&��(69���;��v=�o�ň�`�0�������l���'^�<�}�[�����P�(���4I�G�r���óC	m�lp�4�/r�}].p����hI�y����L�6*%H����`�xݭ�i�F�-��)aQ;�D�X�D{H��~v#����=7�d�Е�y��8�V4��U��Y�ra�>��bu/ue��ۅ}`m�'*#���DV�ݞ��9��{�R�p ���m��B4&)y~��.ٲ�$��� �����}��LQ3k��fQ+d=�v46�IѬkH��E�:�"n�{O��