XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��R�*}IF����$ 5�b^U7�u��g$𲇕�AO��?��4DPo��Y��D�-H�,���ĸd(� .7<�6��T�pH&�*磲(�<*.�D 놨����ō�����ʊ�j�į G�##�M|�`�x�)��K԰9#&���orB����ٛ��PhdA���OT��k��8F=�����7:�g5��߫[�wq�^�c�j��\�CTKg�l�2K@՟@���a��ſWu�"oh�;χ8�I~YRP_�L���~r�6f����ӬA���*�L402�<>m6P�g��M��e��Dl���"��L� �FF���:�;"��It��Z!!�)�!�d�+�c6#]U�2��E�X�z��X��W~j��oan��'3��p~㛫��U==N�w��&ɿ�5��h�9!�HbJGñyh��݂ݞj&�d.��k��/���2DT��܋v��q��=�')����*�N�{O���n���pFr�F��?$��B<�m�󀎨V�(���g3
���������L$d�s�0(`4����n�}�t����(��C_���m^њ?�6��`\�^J��/���C�O�<]�j��4D�F����5�-��=1/�	�6�GG&<1�97p����S��v��_]��r��9��U�����i�HU�Q���\y�o<]P!1��&�L874�����C��������.\�J�v��(|fQQ�gS�}"剺��o�
������%g���+ XlxVHYEB    b229    2170j	�7GhHFx��D�ԥ��ʤZsLqyR�G^On"n��W�@
�ܲ�X����֮��@��LV�2Qԫ�&�1�>�U��Q�ϹT��6�:;�~���3�
!��A��}3�����=-��S_stm�-�K��
ɻ�̯��V�T�"�@�*h��z����d(\�d�6uAo0#!9��@J��h&�|��!�7�Z5X�$�
>t"�����#,?`d�����o�������z��3���]ġ�;����4A��F�
�2$)I���L��\�gٺ����~����fT���B��;N���5�VD�������z�ÆxS� 򖻽ŵQ�W�E��B1�F���4L��s��:m��#���Xs��N@�b�-��#]�a�uF���V�6S�`l ��������?��`W<�������޼/+)2�aZ�,����@�E, ���b��=#�R
�y �Fh��u^p^����a(���<��a+�6�xD��,S!�b�c�����.$�
����phh�s`ɛ*�a*6�S��[t��ej\��tf�V�T4�a�KNI|.��9~���8�DX&�Y[�=v��m�9��� �q�qϒ^��p y�s�޽y�֮��Q��R�S�8OJ���,�x\��������8!x�G=Ȱ������ ޯ�O3�P��迲��@���d�I��k�_�C���7���mI���K��^�K�h� )�n=c	u)y#X̦o�C�d!ԫ�$��O����-�;$�����.����/�ĵ	2������S�yDFB�����WmG!���*�ހ��;a�� �q_m*�8QRq�Gk"���o��	��=������u}N81R_�]w_q�{�*�@r�e�Ђ�#x�uE7#�%&Dn >�����>��+%�v[����-ڹ9k!Bf���]�NCX��������*�qaӧ��
��K�S���m������>��Tt���,=��k��qQ�P���%�2l�7�}e�J\�2vH�F(���LZ�|��Z[���Lh���>�W�)�,nr��NʽvY����s��kF[ϖ/���>�j]��b�����0�3e�R!#�� ��/P��Xlӳ�/?6�Wҳ�l�m�^}���dm��|����w�m�Ϟ�Q��
n�ZJLzcއh��\�M��r.W���Y��{�X,�D��&��F�oL�۟t�8h�1��M����Hl�����R��V^P/ۍ�'n&���n�˜B��ˉ�Gz&nS���P��QB/ƍ81�0�
�V�ta^��0��:zX�����J�aű��R�Y��1Z_y��W�ױL��n���k28�����0)��Y�e�h���������{�X��e��A�՜�}�uK��w���mz9���t�a"���֊�*��as	$�,�ͩ��s����O3�m �Z��bO����mmN�^��Pf���R8��a����q��&Ax��n=h݅�3r�U�˞@�s�@��H)s)�z6�;�y{ilG�<�el�Ȋs��(;0�T�
v+	l��
^��qOh�%:&	��에N�D��6\��*�������u�UȲOL<MGQilK��_'�w�Igܞ*J`��g�S6Yj�K%�0ns�7�>��P���H�Fqٿ���$�ҟ��Y�@7� ����_�C�����>3a8f�c$ҽ����RuWȔ�ݝ)ZQx���z% ���(ĉ��������K�.y���,%3{�kn����)�۶�!%xyg0P�Ֆ�����c5^�����#fk�J}G��0!����/${�v}�����c�l���`:�I�JP�A˓r�̳�`���Ҟ����^��[s�b,�:�w��;f1����(Є�e*8h�k?v�r�?U���[�I�u�����ܿ��Ds�@�e��R��G>��s�o1�<���t��g����|���mk��z��r��ӔN�Uo�^�s3�w��{�)(ʍ��>��D�(6����Ufti;����̀\��E8� 8���"�KB{Ϝ�?��(
���!'���������a����M�3!胤/�hp�od��Ŗ�&@�w�uH�1�&:W�#s�m��'gυ��L3 ����!����<�N�����.@w;�ʾ�ň?wA�e��l�b6�1��lM<���E��c��b�%�bx�0�̜8�c$�B� ��N9��	�3GopP*�� ܱ_�򪮣
��"��R��꧱��Zk�ʦ�!����D����`�8u'�
����h"��AE���|�r3����7%�gō�p |Z��9tږ���I�u��#Zb�ս�U,s�DI?Y'����ِ��`h"pemO}�nX�}�걨L���i�0;u���,136w?Df(����ˊPm�[�?P�V	��=�B�͇u<�cq�i6Ԟ3�aƐ� ���
�o7׺�_[x(,m�醧JrG�Y�ճ�Z�@�55��Qħ��>.�
�{~�R������2=l�m���Nf$RY�>?e�n�7������P��R��L��{4��SuV6�Ds�1R%���[��H��'a2�L�����
<��u���j=�V����ڌp������@�t�m�pEW�p"��͛�{2�.�qP+�o�Ťv�e���k��
ZԏAd�˒ϵbX0�* �w.ˉ9l���0,�:��M	�ͻ�j9�$�H�#S��(�`N�Q6,��R�S�h`���)��چ�`g��ϓ"�``jA>'�d��H.�Ɯ��!bB_�!�~ �(~2c�zm��i�#TS��k0F����¹�l�5�(0��]�O#��8����Eg�x�l�U_���'z P����Ǿ~����ƺu��O��p������}�1\�s���m�"��y �M�i��}B��5YJO���7���m����z1ֹ��Dl�R&�h�Fe��[��Ʌ^�����Es�	��	W��wV�dv�o���6��X�
�}k�`l�� 8宍�'
�k�yŌ�"ޖ`w�A�)����(
���4�{��CT�n��C��2��֢�eӢ�<p�z�+���u�ݩ@�H$}�7/p&4�pk~�M״�F&�=�-y���:���_�(Ժ�u ��;S�]~�ש7�z���Y#�O��P���v�9o[#��d���U`QG���=�Sh>z�%����({�g�܀�ͱTR�����|H(NY�(k��7s����݇G@��<�*�w���no�^��G{b�6��m@\a�����!>!�|���B?���[����.>Z{�q���Թ�.rJI['�;����u��o�ˀ��΂�O4V��`2�{����}��:�Ne� �f�Wz�d�k*��N}����^!����R\�����^���9w5������D�l�mG�%���k����W�.	I�T�+�U�?��*)�}�zJ����_��r跮��]h�S��˗�8<į��FC(����(4���G��V�'����r&�;G,����N�4�i�R�3��vs��Jem�*\qIv�����'Ů|wmDHј��ׄ�iMj�B���zv~�L|��Nd"9�L^���I�����vd�Y"bIy3�M�������Dz����	��ʎ fv:��-�W�r�����e^�ۤ޶�B@�<��هz��֕f�2�� �#����@�y5��U� Vs�I������Aʹr�_W�0���6\j�����m#҆:�%�&S�{E?���	9R�G��Z�"���.�w���Qu��" K�*�ug�����ANQ�t������Hd��"�fm]�#x*3��8���'g36����b#��������g�V�f�g�\cbCme�o�+
nJj͒��3�r�F���n��j��M�c�j���k~�a=n� i�T�\h��A�QK�����v��J
a�%~*�r<�Syo�<�{�|�\�2ºM݅�P���l��3�}�|+��-3�Ӂ�=�$�<^u���g�;u
������ͻ��xJ�ɰ�T��L`��W���Ϋe2��=�~J�1>�?�)&�b���WdCj胊�S?/���#�3���Jޚ�k��A�04+FR2mSy /:�� �n�~���r�Un��O6ᜏQ,U�H	o�[_�D�w��%i<�1 b�	8�x}�MɝGn�B�h���������L�2p%�6�L1�(����rxf!o�x��q7�7'���C�p�2<���n��@�,O_�"��nȫ�V�6J�`v��s�$.#{QR(�׷N;�^y �J3m��D�ϸ2���Bo���wj2��$��K�Nip_
�\!��_�З��O�A�s��L�K���k��}#���TN��ݦӾ�k�IG7(���d�����Q�Uv*~��g"��.VE~K-Q֑z�G�h-߃b�r��cǣ�,7�!��D�=r�	m�?�����Q�ӈ�х^4���P��/�z�*�]oh��"�s�̽Dn��Q��o�+�ͨ+Ws�R>2���rK�GK��x�WϷ:�T-}�gY�r��!�k�1f��4����u��
��G�E�l�-}45b�'�$Mef��?���L�QQ�K|�p	��:�J�Cj'�F<]�by���`��P>���K=�ܲUņ�͚�e� w��vW�x�8DY�k�p���`D�-�Z���������R�V��'O���f��/��,�:����2Y3���>��Y9��Rۜ�2�I1��5^2ikD>P� k��D�@"�Gh��@���~��7�th����,(��EE�(t��}�6���lhˋ϶�],0���Z��A!,��q���s,Sw/p�D֨]d��ĸC+fQ�!t�I�b�I�2.� [;�>	� ��}���ӱ� 1���f�3�j�Փf���SďR� �|�����9YF��O#���z=`��ȶ�����L�ڦ�����y6҉If���p r�u�0�c�GBB�����OIN�z�B��̈́Zd�\L���oɵS�aR��I
z�����]�zשo)�*�_��UdDF��]����_/�t<���<�ɍq�N)Zƞ:!�(�R����E"z�y�!���$�=������;^���}��wŔ�� � ��B�����a7Hz�<���f����3��8֪��Doc��9Ѷ�aG��X��r��Ҍ�!��cr��l����'�'0��U���5��~M��,G����ˆf��.i����ɰ�`�aU�8�QB�N�������\���V@$'U5�6(�`Ald���$V�
�G@_ �|�K����¶F8��\g���*-:A�K�?J�F�E��5�g��)zB'K�,�}L���^�j��CG���4�-y�?��9<0�S�J�����X�(�����U����&[½�|y�˄�q��]|3s��ځ����a�����Z)�X5U����ֲ� eg�7B�fF��|陃~r[��hf:3m�,�~�L_o����'"���$�u��,��������ݗ�a:��HW85��JH�����C�F�F�N���{��69�s��ӵ�e��K��(����a���m]�Z���;d�͢�H���nd�^/���
;��	�b�?�+(�g���t�����#�W��'�{À����cU�՟ِ�[V��O�(-�?_�ϫ �2O�dh��~�S�
����i&kZl�rd:d���_����R9S�ky��˴w�����LIBm��<���r�HGİW���A�H��-q�ů��:}x�����Nx�@R�܌���n�w�C�ͼ�2*��,a��RS��[�/�cQ�&H2Į:�O�}�D�}^���%�������W~I��YvdGZ��4����`���+D�	�ݍ@�@��ΰna��I���N�f�ZKT�w�I��h��3��[#I%��5�t�����>�cT��4�^�37�񷀻W5Ss�Dr#6�z�L*���Z���B�<���d��/�oj�8v)�'���~�1�-�:�Mr��~Z�b�Z���d�^�V�p<y�&�Vj���K.�;Q�
=?��7Yf}������n�L�B�j<g�����łR� �%���hI��EZm��r=(�� Xx�o�ǽ���f�c��Հ=[4[�ݣ���?��&�r_Ռn/e'��	]n�xL~C��{F{� 13`��7��LC����⢾�/dZ�V�F���]����D�ئ�E	�Mo<�����q>�0c�^�Y#�IkvL�3,,
���Y��*w���+�����1����S�"�!_�#���a�K:��TҌ�&�ʴ�7<�h�:�<Q%Y�v$)d��03�U]P��/���{f_�����F<;3Xy0��jo��ԧ���M�09������Ň�.���������s���W��{�}R�<}6!O����D.�����Q���%�4zs��@]����T	Tx5_a�� �\^p����LK�F���P���&�S�u¿Qd�P��?ğTN�)���.��㻥s���tgs��⸽��T�yWO���֖��&<��1�[N��[�-)VFՐ�=Xd# ��&.S�[ٟ4�������9P�n@q�!U���������|��ս�]bP���}��{}���A'�y���G�����+b�|Oɓ�0��A�W�-�fkW��K]�{)EO�0��*h��>
�M�6���]-8L���b�S�F(���L���t�32Ś�9�՛*��k���E�(�O�3�
FX���(���,O$v!NVN�H�t��%��A���ԴU�����1�iicLA�bC�j������|�c���qK�dE���
fI���.6�ksd{q�|��d�p����w��-�H��0ࢼ���B�츱bf�ɛ�6�'2���n�*pA��ǵU{ ]k�~���%�r\���Y�z0l�����	X.+�ePL4Ƅ����}���X�;��c`H�%)����]�����'<�2a��SK����=�
|��Pi�!t����U�¥ I���NXFA�"����B�q��x9ʦ���`�������O��ye��w���mZB�S������|1'���EX�l�f
^
�C,�����x�p��m�8��`�<?��pa����5�q��
$�\d��/?8]E��³�N&�j?Mғ8G�F��}@)����W�[1���~�^��w/DC�5%8�����8!���NUZ����1&]r�@���Ն[6�1��_�Z��]�(�����Vh���P�����s��rͭ+�9�%Y5�[������K(�A�t�A%����e~�_�5��&����p���1��R��gz�K��r�o-8+�{�����/��˿�4�~y�n��wҘ �x���k��D-v�>��(����5�R T�s�(��K�Kل�zh L���l�6O�8��Z
��%�W�A�������K�g� X��ȿ-�z�
�s�]����;��T��w����B��Qcڔ������\kX��[pA݃��%�iRU�����Ѹ�{öP�*3��1�Z'X�^�����T���[�xQ���a�0<sz/�J� ^1gG Qc��A���cX��t?�([Uf@���3�sp�#%�`��#���^����j�\�K��(���P�M�I�"��yN�$buTS�8.m"�8g�/���$X;��#fL���9x�{�*�}P4�.y3]��A�fI����H)dr��(�5�qKg����^w��D6�`	��PyF��qc�OG��2���G�}����H/��s��Ly�+t�3pj��Ӱa��V�i�ǋX�/Dof4i̈�6EkR:��*§�Τ������t%f��R��ה�
Au2b��Kv6?��w�r]�Q��,����Y�ru�Q���d���^.v�L+�g�1�`���A�&M��ʓx�~R��a�el=�#(6��6��|/�@���Fe�A�K����t �yk�O��I�)>7(T�x���� �@b�w��ۇ�u[��oЄ���0ܽ�<�X�`̋H��YI�c�v��W�9dP!�$���D�IP��Q!�+�(H� �h������It�aL���%����;�T�Z�~��u\[��n����=��s�����(���9�b�N0}�s�������|��[�Z�s)��1�l3rn@��F���ԻQL�2_��'�M�k2�+*���ٵz�p)H{���}�^2�%��V7#a5��X�ǁ'����%��?��A���#�(�ё���4�c� ��