XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��t��S!��imԂ�9�D�k?�5l!X�0��ER������G��I�^|����LyGO"��-��V��_�{����t4%���yY�����]���-���Z���X���,.���}�@MT{��܏֙�甧��p�*�����q�-֙7�!��۝��gZ�c�t���)O��8WG�6��� t8P�h�|�T��뷇n�o��|nr����\����CnT���0�S��ϖ�:��a/ݲ9lg��-�{�n���5��Ȍ�b�e6������eT��F�'�`�e q�B�3e�"��*�*�	[eC8�25��O�QiJJteR�c:ݺ	2�X[�@9�v�v�8!t`��}�O��:M�~�Xܖ� �0A����/���gH�QP�s�I��K��3�V��0XG��s�5�[���t���!�u*s6�����\��wf��w�k�ڵ��a�5�s��Цߵ��w��\����9 83n�2������,����},��e|�v�qp�y��W����{�CP��B�} ������J��]�RS�� �"�xo���Ḽ%��}�.��Ӫ��\[�5�vBRfg�]��Fx�r��
"y-���&?{���^9�<H�W�k��T⁤�c�Gk�	}�̷��T�E��j�´ʿ$��{e��0'y[
e"D-�F/���?ﮘ~� ���ͷ�J��-F��-�uG5u �q����l"F�ذ��{~�3��p�I&!1��{�XlxVHYEB    9fc7    1fd0(3}�(LqR5�4�Tخ��`F3�N��YR�6`�^"~4e���Ѭ�{Mmiy�xbយ�ߩ*o@�\���:�t���gy�T�&I.{�{Pa�X-j���ʳ���\fj�K�ڎ�NN���~tZ����#�0��<dF�-:Y�Y�Y+��\�]e���C
�|3Lnpp/��g\��P�9��͑�F���<���D�O�����!�g)(aF]�����0�_������%tY��oɛa?�w�hD4���[�Q=����xOr*��_n��.��6�����r9d���>�aw<�'���m����1���s(�㋢+V��M=.���r��'�/W��{�7�[6�t]�E6p����7�E�hP�/��C���������f��N#=��V��lVR^ћm1���\�U�	BZP�g��ힲ�9����=���֞`yP ��ȋn�m򍇵QƩ�v���U��m&M7!Ə���~���Q�a:�\>�e[�F�)������P[w�H!5��vxL�"���T�8mkS9���`/����k.���[��@rxq���Zt�����W8��J����D�w|��o�&��s�p��6���^��ޢg�_آ��V6@iX*�^).N�
��pB;�d��N�_q�XE���^�
[hvP���l3���vJ�����è~͖����8�~�~��xͽV��~ژ���h:u� }��k�(�՛�*(��-�	0��=�X����.���Y*E���~�9�,�����֌��bϢ�R�B^%�����Z�v�1�(6_�`�	Ω��`�SX�U�P�tCE�|�=����)f��O~`��%��������C!`m ��?Mas	�[	��}qF�VR��7l�pM��\k�n�W����
udƞ�u��,a���җ�g|	�H�'�e*�_�z<~1�}�df�tk�k��ձ�Vn~R�x̙���x@��>Ҵ ;��%�WR-���\
��8#$�����V[2�i#}zPNm!	�1�ȫ��N={���c��5����.��⸟$�Em��!�k����~~��<nSY~�W�ֺi>V�NƋ�;��a�w���)<@���������[���[N��O�q�q��G��;�"r1Ϲ���D��'aĪ#���'8ͳ�$�h���RmC׍�W��?�nʅ��3�c�L��`�_�����*�j ]�؄S�������&�o@��i�6�./W�n7>tcG�-2��)�t1���w;���3n�
��t8�u�� Цw�;��Z9�ѣ��e�e<��"Z.�����E�B��a���Q����r��#b:Ќ���l{�Ɗ��w�yK���IА&Ym����?�C��΋�?1_?�hY)qu*��A��"���}Y�i�i���|�L�_����3�)zUc7��X�`���D&O���=&*���!��$��D:�!n�g)�[F-�Ǫ`���OD��E��6)��3�y�ȱ�f�5�0�x���Gnʚ�M50�o��>��K
/�\���EF�Z<+�%���q�V�G���/�1rCubX�	�
������W�h�̃���dҔ,�,��n�[�_��O�cډՓ� �)�ĳ��ׯd�PK�NK������T��C�w�ݧ#Ǝ ���!�N�Olk�8��pN?�E��@ F��	,U0g�$tə���UfN�x��1��W�Ő4�D���Aݪ��J�/�?�˝�"'3رG���)$u��S4^/�b"}]�ϳ_ȸ� j|���+R����J�~���#� ��v�!�%3OC�4�a28�;��k���
>�󲭻i��;pE�:�>��v�Pu�m�������;��zS݄\��\#muo�z9e�ԛĐv&��џf�� [6��K�7)�N�"���p�"��x�m����$in{ކkђ/��v&F�h��;�*���,�j���� 'e3�p�79IJ�c5L;��\w�|�8d��V��A.%�[�lB���W���<);n�<�eW�ӿSG�7jݍk!D<�w���:Nf6�*F&A��Ū��d��E���f�;��[I�� �oH�{+��oB�.�q�����,(� ��E�y�ݳ��W����B7*��`�q�W��@��'�jΈQ�@ҟ�e�? _��U�nmaD~�fGe�%$5��-��'J�������Z����ŮjÌ 4z;�쐲�.:� ��9�M�B�Z
�i��p��`.*�9���g��ɼ�J��� �*u����7�i�}܄4G�A$��Q�����b�)�cɌX����\��^1���WYV�mϡ��wN�Z%/`OA��_�IW�~#r��4�!�
��V\ç�u���|���� ���,����`��g�2����\bʦȸ�U|�7�@�������9W"�>u���֑���Tɋ/W*��<�$��n�7�w�U/���µj���s=+�/4m�	*`؟�;�O�Wğ^fOP"�Q��s������^z��0��CV�ƵYT{?�B�gR.���u��3+ɨP�����r����w�"w�^�Y1������3�C_����F+=�e:$ӝ8@�by%���%ND��B��'���˘h�ʩ�����`�%,{²��0+)oom�#C^-K�m�_@�U�o�-�j������9��?v��P�F=��ov2@u7ь$�rW�TE}��:��P��IXQ��L�=ߓ�3�ѡ5;z�L�_q�~�!�]�x*��5&~��?��k�UԄ��h�`���`!V�;9y3�=�5���i4�b�	48
�ή�k>��&A��R�\�{	mw���������{�1q��ǹ�6R?	7s�4�[���쒓�˙]g�q���+v�7��Ӓ��,����/%���?Gh����px&�T�+�N�D�󹘦����3m�/���eV'��ͅR[��}�GA�����G;�h��-��@��xO哖�M���:)m%l��R������+�� O ND���T��� �,�7�y`/����u��"OQ"����̨�q�7�s����+�n"ā�/穇���Cd�8���>>�H��Se����(�r�\}Z�~���ܡ_ax��|�# �ns�<.�R��w?ꧤ���]�H�M6���&�/�3ȥ��� է��c,OuT�܎+`�(<O���Kүv�����c�� ��"��'%��~��3!y�l68����k���:��#Y�CXm
�)~HΖb{��(�W�y|�F��zV��ػ����d�̺�E1�W����A�����]jq��w��x_���N�������oK��B�/z2��i'��.�)��b�,S�����Q��԰T5��!_+� �A�gޮ��	:+LKz�.���
=64A�)C�A��`�=�S��~�0���L9�I
��߹�-QHO�c@�S>�$�4�}[��-P�G�g;�]eܡ�(�-�r:W�Mb����+�.�a��u���2$D�e�y�.����⾯���p�礄�Q�0x�V;s`-�b>�I{%�|n��㒮�	��(K��8�Q5�9�������Ӣ��\X��s˙�u�ɾFu].R�}�<�в(�f�Ւ�4ޯ��M4R�%n����6ï>h��-_� Qn�Yߨ]	��,7�g���bf|���q���L%����݅�����;
��H%��|,"���^0�M�Ź7���,��B�,h���jTI����i]������Z�e��a��O�BX���z%��6�i�0���3fQ�ʥA���T[�#5����	��� �s���$�z>q��0��,��������Z�n����j�Y`�6�G���}�
�{l&k�S'�ޖǈ��9�N�ٴ�jܿ�1c���i���n*�BD��]����i`�zHD�j���z"�(�������'����#�����P�EJ���uw߹�z���i���r��!�I�j5�-%�_���N�_חPV�~��;aN��'�ᑧ��"2��_�I�A^#��E6�q�ձ?6İ4$� �Q�*9��8��$}~z��=֐Q;\��(|3�ئ�c�r6�/waV�u�W)�#�Q�|�o�8�Ѷw��ﳹ�6��̐�٠W�|������ȴM&z���)(�$�N���u<%c�DRQ��[���!�|�w�b����݂{�2��M��׹���F����᫟����xwZ8��`�4�A�����m]a�q�٩�p��AIk��D������*�%��2��~���\�����_���jÉo�B'��A���e�OĜ�+p&����x]	�r�ݐ�������:xC*���c+p��b���
�"u7�s���o8��9��s��ѥ��U!(���;5��7?�.猿Y�sW��SjrE�+
�/�t��Kc�]��ϺF�t��pN��!�l��d3�AtmD�z�1~0]��&k3mQe�ڋ��CR��S3(<��x�'{�A��XMh�b&xh��bh��K_�EB�ב��"�D����Nd���:��a΋��d�c��}=0N_�ɕ�r)���?F�2%�(Y�L+h�@WRKsu!T�;��'�EKlDE<�2ص��wҵ�It�0�Yo�7F-�p�Qw�����8����T�4xa�{��6�PEk�6�DO1t�<�����J��r3n�E���5֣4Z��ۡ"0E�	����	0�������� F�>��~����P����IT�#���I:%��e�¹{� ����AtW��ki�$��	��j_��|D9�����i�L��\(DdUL���:��i�P=D�\u�5<D��P�n�|���]
�坁&T���-�^~>�:�l��ȴ�X���mAT����u���}�bPI��y^��סN�G�X���ܒ�>�P!��3H�=B���1��&���*I�m ���s�oX88�D3ZE�� �t+%4���BG�wCb_�L�P�}�
`:��
��@��g�g[��v!B��yD]�X�������hƭuڅo�A/��9۬w����7%e��lR��j{�6&�:Ja� Z䚀�;G�2[�#����&�-d��=ڗ~P�,� Q!�%��<�%!6�C9��/ߎ��+Tx\5����,�G?�հG8c���U�j���/!��E���10��)L-��L�l�\	��r�$����6�W �!�؀�SM+����O�U:xW��T���.��Y{�-.�,����#
~�A@�.h;`(��~�u�@�C�:�g���`�]�*V�d��I/]�~��������
�پE+ș�-u���!=���:� ����i�y�Vj2T+�$o�F^Wޜ+Go.�jc��rژ��/�E�;,�F�ݑ�q�|��'q�^�*G���J�=gb5U�Y�WM|�S�����j�ե�0��@ΗZ���`Cgom}�:�t�X4�������Y���pϽ����S��?�]�s9�b8M;�-����ZW.�֦����U�;YS�N����+�4�f&��t���a��%���6,�g҉d�����B���0�O���'\۾03EkF�)�iz]��y�B���:L�̰�FH�6��I����G@�=�j"U �'<K��Ŋ`���g^����ਇ��L����o%T��e��0G���S��(j���e�&���|�]�����OɴI����$H�^��ڈNun^�a�� z�>O�s1[�N�}M�^�(�1�F���$B�_HR�q�@��k^pȗ*��L��K�M�$��dXj� �[�,�xQ���gV,����~�:'�;j`bV5T�*Ek��kZ�*�3+�$k3����*��l��7�B0�6EK��߈���{����$��#|�?+�J"�y�~�-���G��Y�vD�v�^ɓ�G��ߍ�h�\�_OJ����Pd̼'��}�%���0��{x������]�Y�Jx^�X�$e^����Ip��,<� �AvA���MH>�<5ȉ`r���C�~\G��2H{(���*Fh�:���|_���6-\p[�v��Q�/\�
zUYD��]�f@�5���RɥPZ��U������;�g �"aW�u��D�֥������4O$?����A��֯�g� ��:��z	l�-s	��"��=ԓ���(��(�K,�ʳ�W�����8�����r�l��p�$<�g!G�>�&fJ�xjd��C�
u�h��}�O8���e��\�δ�9���h�{/RJO��6W���2��̎�b_	�f�pX?r#	#7�Gf=��p��x��,�����N��q���$�P�(���?Q�+�!��S���H����9��c��9!;(*��Vf���u:��Ӭ��q�7� gf�y��*����Z���x:�~�D�]p�+�̚�f!���CZX�2�T#G9�Q�z�S�����o8C� L;���p�SVa�%����4+,�b�ϣs'��d"�uAg��������f�N%!�:�����R��LZ����$bs^��Ak��9����x,)��aSQ���幼Y��_�a��V'`�6`A"u�gy夠�M��ۏQ�Φ���Ah8�>Kvm���1�_�,j$�9�k3~_���e��́��=ڬ�U��{��� ��_:�s~f�2�p|x�����}oP����b;R�Ym��#$���'Aj�1�?!�5�vH=��Q��*ҧ�ؚ&7��M�0�\�BIȩ��66�۲R�U�t��]
"���f��b�:��溆���c�v�]2��y�w�s�jH1=�R$Vj���FrS֣��E:�b~=9vX5/��/��h�䇋�t{=�!_�u���ڎi��̫lΆk��(k�1�q٨Rw�}}��Ӛ��N�ίax���j9*_�N�#\$+���~��p�U����91�ǯ�.w^7y�;���`�辗��u,8h�#�r�����Jw}�����_�1��<H@$	}u9�;�1��`��������~�X�./ڢ�	*�݊���Uv&��2�<��s��-�d$<Fnt�0m��o�BHM�*K�l�>v'R�Wq�K)!s�G�ٚ�S���9j;��]�{ۥF�>��F�� 3��ݗ��*�X�}{��]�����:K��Z�� _ń|��q��.�Ww��L����?��uŝL����,E$�I�8���1�ɦhҒ���#����N��+�ۜ�O@F�H�dΘ��)�2y���i���l�-�@j�yT��#��.�d@�-sK������HL������Mj9��{�#
�/�q�[z��c��b�p���]��<��{'�}B�@E��=�9ѭH��V%3�;���e�H_b(�`�Sb�� �~^��Ѥ�2'}o�d�C7S�W�Y'�Rm���e��4�o����p�3���<^�&���$�)��\M�NS�������1�qJc��1���$�,���%()�!�щ�qID�Ob/=7l��`�`n
����U;�/;��|Y3J�V>�)��Zym�Ǥ��j�x�� 4��R�����Z둉��6	�4��~����N�l��H�$l���$����ړK��ګ�[���}^�g2��8��#�;jdi	�B�ܱb	G����[֓��P^w��1Ȍ\�i0XC���z�v�(6X3�$��D�'s�Ml����= �CS3/K�^ �_�Z�x�Zs��]i��$�:�X:��B�6�ϸ�����I��8N�X�	U�6a����P_R5jC��d�-�~��KҢ4yo?�`�
�1�Em���n=�k={�Z+���]'��`��c%3��P�.��q��v���T�����k4�oM�)�˓'����iw�-��`�|��v��P�s������SyJ?�C�A�
�툭��� �w�x�U-�I��脳�����n��E�m5�_d@yJ,���Å��py;�"�0�&W(��-