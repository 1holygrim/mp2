XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��'������?��]�a���ug�}5��~Q_��=w�C���-�S�����(ŷ ?W�o��x��C�hn6��d?�I.��Pc4M�Ջ��_���L�gF�f|�F���g����~�*�� D���٦1p^�+I"\������9೪[�	��R�a0�V��Ҟ_u�X��e����ȷV�X���>i:^���	׵k��F��s�\���%��Z'?H�Y*\7���Mcu`��0@qpя���_V0��0��YO���9Ԫ��W�H��\�k`5�i% ���0u�t��>�L5��R��!�L�te��.U�u����F0�y��X�Y�з#�Se��S�����t��Lخ��d9��I�[ʻ�_�!݀��Je�v�#���t��apu����2�'z�����zI��K�Ě�C?�L��~X��7�sY�vQ���%���l�b�3��u�r������>Ͱ�d�i1��/
K_�i�6!R����ej���־�EJb�}\<�w��$���j�x�.έemI�[���~�1`N���<�3_����������;��k�W�B��c� w�e^�1��z��i���f]��(�-]�\����xl��?�/�E9�b8��3�8�ʀQˆ�{�,���S�y�DQ&�,�^j�q5l��K�#���EȬ7��S@4�D��ɗ�O��m�?�b�`"� ��/��o��!��nՌ�W�8�ޯ��K�KwJ��f2Z
����?mcXlxVHYEB    3fdc    1160S2�(�w<=�qj�����A�Lg��u��Z��ȹ�p7�[���({���O�	;Νީh�6t�P�ߌ �v���	�>�'�ܤ�3�A����ùB�(iA�3#��c诏�ʗk:[�g���P���R>G��N���#��4�jC�}J����m���̞{|~r��p��9�I^g�̅Ym={uCz_�2hL����4k��$)p$�Qjn�]|p0QY�"wg9#ĺ�m
c[qƳ�J�|;�U\	3�C:?�s���@ �c�r�7P���eaB�ɳ%A����t�k7)�!N�e��~��s�R�hM�>��bp����ŗ�J���m�`(Z�p&��pv>hc���<��B�k=�r?p�H&��FЉ���ٷ��J��ϔ+�98�1���ژ`i,���aQ[��R���?3�j����৵��T�����0$��L��r�Tm[����W4��H�͋'��+2$�"�yX}bf�n!��T�������X����f�]���sʳ���N�]��ؖ�L`&��LdjN�(��]W���.D��Ħ���ͥ����{uma�Z����ԏ2��T2���]�r�>�h���֎�Ep�(Q'�Ȭ��n�z��`�� (a��V'|)+���92Pc�n�X�i���=�"R�G�N�������{����۫��������"���+H��L�g��wFF��篙�׼��{fT�:�g�j�%[o�1��̧�1l�����Ԯ�p}S3�[�Gy5+�a��v���JBw!+j(:�IP&6�2X��B �zj,�]-b"��ށ��F���-�U	~�����%4ӑOESE6���RKh;����rʒxSNԀ���#�f�f��.x���s��S&�p\CEϭ��I�°�Z��<�t@�}�lO�i����30�+�e1�.)��C*8��V�s���g��]�?t�߿�U��� e�����P���������@h������3���
}���^����'��;]���p�	����m���}���sl)Ͽ;���{�?���oz=��VaR��"W͆�7�5y�~�w���;����#�{՘x�~;H �1��S�u�Z�x���ͭ�o�ʢ�e?��=��~Kf�Z#��S�g"�\.��9�J�@�E>��{Y�C��V�,�]���uB�z
��3�n�$ 5��Mǂ�����/���#&d=�.���So����دdC�Z�H'���vj��b���c'��Pt��,��+έ벲=-N宂{���0�V��G���gE��E�>�{0���Ǹ�)P����<%:�p�W��k�|��c��:>D����S2-�q��M$�^��D��Ӄ�N[��i���`92���	w�h-�ф��H�ͅ��r%w\��&�pStU���������V��f������X��ʷYx�ob�SΘEg��|;����:�<��?otcl2T��u$B���a#_�?%<�jP���Bu8�z@��@�M�|1�t���V.6#b_B(f@`I��(�T�,���<�e�㻭��g�r�G�A?��?�r�+��s�v�_�����b���Vi�,�5�wL��(�i����a�ZY�gJ��s�4C���Y�kY�N�Sp���fG�e��".fu�� ��9E��'�c����K-��y�a�>��PLK��1��Q��d��_�<6�=^��IZex�x�藤(د��X� ��)�Q�*�7���oG���'��+�S@LL���J��Xh	�ɬ���|#�&��(��ߠ��_W/bfr7$>��T~¬��7���?O��1�~�*�Y�j.�W-:w({�	j�3w�B�=��t��uy&�w&:c�7�A�]Vz��-&.��h� g�*P��޹7 ���a�hⓞ�o�܁� 볥��w؎�� ����m�0�`Lp0!�Q_&�V6 �P�ʾ�+r���$���>T<�]�JE)�a�m���#�j�l�Sӥn�⤨�O�h�?%�q�E��e׉xQp'��r����J�DYdC�򚏉1B��a�G���N��0p�tM܆Q	��?7kO�CW��.���!�ɘ�x6����˺W?���e�x�k��>9��Z��ş�z��Vϡ�N:�1���xIJ��]u�rV�C�a����w�]�R��R���c'��@ P/��+�%w8l�V]�{ra,�'�[�����m�iJŃä-N�zf%��q�u�m���;%c)�xf�k�Qu���fޔ,��:��e�����e>g�o�5�4 x�G7ꋋ�nW�,�e.˩�:��c�K%�()�h�+��%Kι(U����a 5��z��x�)WtW�~� m�s���$�[�N�7HF����&c�9cєė�g����Y�W�[�5��}xfn44�m��OSg)�mv����D��r�����d�g��G���=V�x��ق@�D���w��	���� 
`�
�{�ڃXS�\O�y�%��[��|��o��6�r�|�>#���Y�^�J�R���Hdx��{'�WI����t1WKJ��>�De����C��$	�(�&+@�r>�c�ឿ�ő&o�NDb��;�J���6�|�M�� �}���h������i�=L�`��G�9d���4)&�.���h[(��Z��<�X�臕ņ.ܢ\\\�]��v�Q��Ca Xj�%��0�)�ի�r�1צұ���Ol4�e�S�V��~��d`$��xs�4u`DzS5�o���- �*O�"�P���Q?������D%��&d�0э\�C����V�੔�0%��i�����X"�p�yH���Bu1�K���:�U^��O���c���f��t�T���.�di}Dw���� �%�
/nڵ�`9����a�2�}UME��3�Ⱗւ���I�C�ߥ/7*fh���8B�v�i���R��چ��%|Od�㓀6������+�Fn�����F�z.O���I,�X"�H/���P�<�#�h"���|�:�N��N�.���LB��0c_0�o��$�Z���Ho�y�:���K�C� j���S��MZ��B���a��Z�2�$���pyE�d�$�zo|����kE�GO
���̕t�Q�D?_;rq7�i����/B�e(���'3�g�n�$��xI.��݇��f������XF+���,ϝ�6����j�dWb:�*��?�K_���j�'/�@�I��oG�bQ	{}���)��*�9�?G���6_�ig5Uf�u�`9Q��Ɂ��{������R�����B�M�@�!g����Ӟ*o��y�,l��������yPT&��9`�d�{�Ѻi@�{�)K̙� NC���w9ۯ��S僽�oh'��8%��qYN�?�9c{T/dmz�S;�T�"~�z�H(wޫ�V����#�K6�[�ŷ]�5���Mz&Z�M��!"���V������]�Ts�+����A�4���_G�^G���9��,1��i��D��ŕF:���&��Y2w�e��}t�]����3�"�}��I�X`�ԡ��M�"��O:,�Z�uׯ����/������e�H�h�G*�����8�a%���� �w������� �M�$��q�t�W��(̞��f��s@Wjf�-��S/o>J9 .J�?X�B�ZV���f�6.6^�8eM��
�mUL��'�0lJ�9��o�n�_}E��Њ�+��H���	�Χ���Y,�np�Jh�h�x d�gl�n��X����ߜ���1p���(��D�"�"b;^⸜'���f�B� m�̜��ݛ��Ƽd�¹q֡�S�ǽQ���X�ݪ)b��Y�6�y���R��ZN��V�s��pV�p���	�ݣ:�-`�p['p`��*��Eq�#4d��� n�e*հ��}$s�ƉjF�g�:�4s�X�)bdr��F�~8�-����q�u�pMR���u�0G7r� z���p�ZH�����,%�'���K�������R� &�1���)+�q?ɴ�����6g���Y�C�mݙ�x1�g1�$�s2nYz4/^&������R����f��wk}y��Ѧ��4��o��C`5��+6�7Ī���.iʣV�鵵<NV�ڲ��\S���A�8>W���ⴍ��JX=��k6fGXx$��KQ�����wC���[t[��t�,�0>b�-D���3�7�sە��c4*�.�}69J4ͧlh�����#�;#p'��g6|��Q�	O�P��!�?��%o�h1g���z��.V����<>��L��C�8���Tg�h�G��QR��@��T��X��g��6���Fn����