XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���JYʬ�9�{���/>Ԛ\ϸY�����(��0},6[s�0~�����&�if�\�M�'��w?g/�L.s���_̱t����Ҫ�D7A����:�7���<L�����ϠI�k�ʊ��w��sUIM�Zi$��3�ѐ�*���
���'^����O%����G��(D�Qi[͹���zL��L!�eIˎXj����*��=�,1�����m��F�AD�)@i��mi��-{u
���l�&U�ƪ���瀗��^-а �´�h澉���}o.�B5Qf;���d��G�z�g�6��NE]_g�þ�D��f&��"�T('j�k�/���\�b���x@�Uq\����uIQ���N����!�g�k��~������g?���DV� �Y���}�c�Ju��y%䏨4�k��Wf�����ǲ��Es8����3���^a�I�
$��8��smI
O�B�@)�0cQ��و�k�E"gj��>/�B]K ���]�X�T���~p���K�	���������z|���DŽ^1=��rn��y2��&��|�_[M�9��	i�|&�'rz�w���H0�|��� h�^ENA��X,�=�4{���vi>@sGf��D�DF3hW���P?'6��w�����G�����֗]�u�2�4���4���h}��$u�/y��o��MWy�3�E���KHD�7��P�B ��ɩz Х�tMIqM�%S���`�(�jl%�+���</,���v���AH�XlxVHYEB    da59    2e30�w�����{��P������%+��[�[d�P5�%�"��Q���v�^z��܊��0�VL��ش�w�����%��N�QǷvM���-��iQ��[�SN��c#���A���Ka&%�]����0�)=�s�JXό�,�R�}U��S�:܄��y�\�|_fs�> ����� j���M)@� ��2��"`0)Ao�'/����{'+e��`e �ۤ*'@d�"��&N������b�d�Ln���MY�ZW��4ZlԊl����8>��������cf��M5'���bS�e)<--u����˩ib���Ż�X&�䰇�kf�|,��i��O��ee���#ď�޶�,��/��[6�N_��(�Z�&/�4S��ۘ���j�ep@.�	�#����Ζ�٘GK;4|i�3�2���CY`W�J����m����g�+���8»�i�!�2��l���N�F�S��p���6NA�SmPa�w�R���_�)�.�2��8y�X��x�@OR�����2��ː)"{'(|>k�y.f�(r�ю��bR�x���3gݎ�~\z�f�ˢ��;��cü'��,��fd��k�$�����7���g�h6W��0%Is�F�����~'"?�!�#����[�t�ʎNi�������=�;:��M�Pe�멀m�(��G�k\���͓�-1�$6��U���ɨ=����y�G�8�F0~:�I=��&����(�������g �I��<�	�)D�j�Oі��m�@겕�0-Eu�����+�����q�3t��H�
/?��Q���/E���9�� X��9:>�����Z�	L 	RB]8��KϹ 4qH������\������ƣV++lIM��hz
��uZН'�V�v	��ۖ��<7>�DTH*��	�����h��� ���_%��C-	q�@�N�+^�x�4!n:*�k� ����ͧ�Qힼ"��L��b��ş��L)�-P!Y����$$�l�q�p��9���%0���n�!ԹT�6j�lɗ)��gl�Z�5�T��&}ݶ�@��6PY�ţ�*V��M�>��C�E�-����V�g'�k#��:2h���/��LP<�|�kCy���yg�C�" D��߱hoo@�kW2q����Qe�����#��g����A�sA�mj��o{�P����u�u��l��\���vQG�Șz`r�ު�V��:'�|.�\���$����J�������l�$&�Gn�lfz���g����y�5�d;���/��RY�@1f���Sܧh�w��8�oRN	��N��?C'�]�L��>�&���W��9���EC��b�U�T�z ��P,��HS�^nq��|kc扚�gP6>��\��$���K ͙4
���=ՠ�/��q���-��u7��%�_�Α泊{��H����L2��hm3��7}�v����p[�#�kKuT�B�8������ڎ���������p��;�<���Ki$��~V�R�>Ӿ2���yfE,�9�Z�w�W>����~�dA�0��;�0���~
p�_8�۷R$�$�,����U�L�ե�k
�&�PC��E���s�<����{p���d�Dg�{8����߭'�\S��3�o�������S�Do�'	����ꔖ����7�.꜅��|���6x���M,h�x�����*�K7�ԃ��rN�tk�����.s���v/]6[���2dd�Q���M"�;챈N�Ge����:(U	?%>���W�BKP\��k��H,;�W�i��tI�Lُ}���N���V�}�ql��n����a1�l�N4��Fw[� aʷ��\��-��s��p��hK�A��QDy�c/Yd��h�4�(�`��QFγ�Bc� |�YԗNڽ�E2Ӡg���
�UP��$�j�s�E�@ ��j06�21mܭ���yt��x�\��>>E�@��57��u�cG��R`�>eiA+߄������~��G�&
�9ްf�\}|Y'���իܴe�"\�PF����� +�ȯq
8��n]֜�,����2T�~�������ш��̹����`�4�XW�E�����V*W@!�R���7��N?��~~轔�Wޝ�g�����8rQ��u�ר+�aZC�M���ݯz��-������-�V��N���w;��z�ZZ83�_���AU���{-}�f�VPO�׈+V�>O�j�9%]V|�!�$�z�����.m� �&\p}��LHI.4�U�J`;���W��n8��2O�7됎�F��$�Ţ�``}J5��� ƱN
a�䨍`�G,��Ӌ%�g�)3o@�м�;]��h*�J�Bxk��9/y�,y�-�
-N����I|C����BBɸ�]���s��&��<_�j�9�ڏA"S=�����0(e���3�IA��̤��k�?�z����ڃ8_�d�p�wx�U]be�We�<>a�����KseR������0*��4��y����&q�͆r�o��]��M΍��W�#�ye�`ϼ+3.S`���/g��
t�j�	�]Z��N���xxٌ��ޗ��������i�'�{:�e�u��U?�cή>��ʔr	G��"�� �UB����|�r�E�	x?��GD5���t��P17�M�R-��O�_I�A��jU�U#����~čm/���Х�&`s�p��nUR�	p_)�G���m�I���$���cyἡk`q�$�>��?3�p����h��|%�՟'��������|yO�}YW2[{�mu��c����صpҪ\�����bf��C9��`R�k�L:��,s��C>e�y9������m�db{� ��k**/�خ۬��L����L�A~�����L?&X
��ϛ�`���O�$�do��!�P18�g��rްc=mt_�%5�}�	��*kj�/�5��T|�Q�g��7����jÊ{��"#�h��m�� �-wl�S~�2Ɩ���.�.D�1Ϡe���!�懳���v� b똩�9L筫�}:��>�W���~�<:ZI-��57���"�cQ�-T����F���	��)aJ�F�%|���G�u�
��2��]����<�R1.�5���Ƥ��p9V^������ߔ݇�v��\~�h�Ni7y�<l;0��vi������1�}L��nʔ��X��Z�k���7���i�II%~+B�)o��U�uPf��[�Ec��bsA}T��E|ʟ�g���f�YE����N����S#��e��$�0���F���;�Y�L[���3:�rƫ�cbC�������U�1����&M���xj���hH�q���Ij��0���vi�v4����vC�Fy���\`�OTa�u-Xm4�}%DW��[rJ����y�M�2�@��9�v������39����?��U�ȳ�MI&녑�����Z;��)L�~R��/���I��-��<3��ͣm�Ca�b�c�]�p�"��5�Ԕy�P�;������A��N����s�Z�z��BoWWm�U*���54�y��^3QÚe%��,P���
�\v=�tS
���h��f��a���"��:21n٨��o�	M�+4��F��AcF�$�Ҥ��zq�:l�V�o	��''&������Z�$2�{{�� � ���P�% ��R[z�N�%\�
��g����#Z�R'=���鱹�r��Ғiq��Q��J(Iv#��$%��̄z�bc.��:Q9~	x�m�\=�1'�V:L��r[��G�B'�Gx���J"�w�h]-:<�-uk.���mT��=X���Ew�>�:�����+�{:E[E�˽�rM��	k~'�]U��iRŁ�t������c�k�d�"�!�')�>����M�c΄p��T��CH�Wv�b�qן����'=O,�h���]��hu�2c4_Z|����h�n�3�y10����m��	��j��٠@d/	i��*�Y��'�d����ۦ�,����P��T�k��zC �`��3oz2�	����4l�rp�'epì���$�O{KϒX�{՜��4ml����I�Td0����j87� $����|]ì��cfՌ���x����D�]LD
�Z�F���m�l{����<� �e�C���[�_��w����»���_ �˪�� ����tU��B!�|A����Ý����T�vc!��۹�F��eИ�"�-�T�q�eke�l���M ��Jf�����'a��0�n�67�yg~��Tu�R�3�9f6$N72���CcQ@$�r5���Hm�ĠNg���g�ZS-�c�A-x������@&RS�($��b��m�莫�V�7J�ǈ7B��K��݊�#)
ۘ[�J7,��I�]߄<�' �LLÂ!�Mk�R�.���*0P���f4��6S��[e5b�D\����G�y��t���
5��v���8�T��`�s���,���װ�M��*�r�5��i��'}\�u��SH�Z�.1쾓��.HcIT�V�����נt�Z>�0�l��TM���נ�CGrow��l�,"K�SX���)~�1�&QPd3y�b^(����������y*:Z]ƫ�@�g����:9�� <��6�}�u7���5��Գ\2���wM
t�r��=� Zn��T�l0����MU�+2B��?�O�˅�{E�y��r�����%'d~�ٔs��+v��\�6qUU�����o��a����x�ZS� �yP0�ᜬ*$V2����n;�'���XW]�3�����x(G]8���#�*Lb�k�r~}�{*|ǐ�,�9Q�����9�z�3�=S�Q2�����WҼ�<:�!�����["��M�(�`b-�c��h�da���,`��){R	�ď73\�A��!I���?�WM�H]�&��R�:�\��PWQ����ړ;"���&?o�n�/�u߳������6Jv=���m�cC������$;ԏt���u�� �_�OGq���E�ߴ�O���1���0�q���rx|W;n�
��	rP���~q��n��k�XY Q����r���*�p"Q���E�d��蠽T?:��W1�ٵ�K|:8�(=i{�� ��9�"�q�|�ύ{��Q�M[�����3O=��A�t!?�	3�~����t� ���0��"�k���_l�����h� �#=�a�mr֍Z�E��p�b�1��&m*�WnQG�`�E�H��,����-�	�r�S�w����Nځ1����d�X��������~v |��I���ףz��,�s�ֵxW^��={�yF�fx	����F�/'��#{uM�Nh��DA�D�':by���X1-zb��M\�\b��ho!U�sN�c�Ip�t��x�� h�+q��V!J0����0�w��C�=�aG�M+$��V���l�t8���Z&\����O��Z�CE�j3�b��ivj�.���?�.����
��؉��4K �J�X�0CʣN�&��{��$6t�Ƴ�RJ�H��3������mT��ٍS�/�ʞ���.��i�+n�k��a�/Xjt���2�JV�d�%�=:���%��STk�N1�_�a�p��¬]����h�m�Y��!�a���Fy�+1�s�4~/�+�{�l�1hǹ�&���o8�0}�O�) s;�E�fFfY�Qa��9>��������Y
�W��m}S�Y�̔/�a
3`�{nJ� ~g�H�D�S@��٠�4_#����$�K
(�@��X�E�C HޗG�U�����Ւ_џ�7��52oD}�_�m`�Eè=�X"��M'f��&t����t$�W���yc�Kк�����gS��R���X�}8$O`�C�rgAM��҇���6ɼH ������)Kb��%��:�.��t�d���F�jFn a>BQ�ܝ惝�%LiWgMg�Vo�n܋���4�Oj��we@BUeW��	�\�\aՌ���1c.`�%`�_�m ���#Ο�gq�J���F]G�g�Z�䵠�����5F�����,Ij�)-q�����ݞ�\��H�.}���ݒb27�A!��p��jO�O�v�y��&3�:,T�����,++�W�rY]�X���'�'���"u�A�]P�
�U���,x�>�O��������zg�mT����p2s�1�P �����?!Ͼx�������Cp�)�m罁1��C�-���٬�dt�P���$�Xc����o��d-T[���:S�o���P\�( ��;%�:Xvn��X�Z�I�orw]\Ɣa,c�N��e@���D�����\����G}?�W4���]�tPW.���&F,�gg�rq�&^��w�4��׋m���{r�hY�"�	pW+��z���I�s<;�ħc��$��$;�Ő�ޖ�3�Ma?B�
��"�{=��$f-�3���Z�x���e;v3�U��kW�β���vG������:=���ke��n����f¯�~�/��+�>����}��4a��7 {O���Y�\i��kBH"0Dj�I��'���!=�z�A"����z��H,��`���5�w�\⋪��p�HZ�YL�84�xH8����Թ�Ыz����Y�(w
��Dx	*�	����(�����)�����n�PUr���D�U�k�R�Ȗw%2�F��M[��89 O��_=�ސB|����v��Hs�>E��e6`4����P;�o�͛~��p�<�(\'W�~���ZQ2	�`�tA"�ܘ6�n��+�B�(��X��`Dс�9���S�+��2��M�1�j��qk���2r�<%Dq�M�o�ĊY�G0MN6஦���s��4�f�+�U�+O�<�J�_k�D7��U�wL@�]�*�
c3���@ JBH��Lzk�-*U2��<# �]Al?#�-H2։�lRWz��[�K_��=��PG�-z(&� ��mp�|HD�kr9xP��ّ��Ќ�7F��0��~=k.P�s}*Q0)�����Ʃ����%|.�*���W�a��r~����j�TK�v�W�JS(�:f7�0����ƥ?�۠߼]������}���eJ��Q`Ui7��|ێ۵��L��0�4½y�A r�Ǟ'f����Cʂ�\å�e) �H@$]Vؼ1@���_No:��M���'��9x��"�����$:�$an����Ұ���F<wn�����%pl#}�P�b���O�A��Sy���{�Ղ����E	$�6AWÇt��K��ի�)[�����w�!>T����\"М/T�S>�z�Vt���DV�_~�S^��]x��=�e�}β�kga "�A��_��Y�@R�p��Y�8c�(q���eJ�=��B����&������!v{I�n�C������H��jۡ��S4��o��H��g���O�C�Uد�7
*�y;ʹ��oc=�آO�J�)����1C���V6�܈�f�:ϴ���o�G���%\��=q��M~\t���X�`Q�ew�Ry����!�(}�V��x�($q0�?��1� h>���X3߰�+��U�姿+'��\�Q�����%O��2��l��2� ��<��Y<���U�ܸy\4�����H�o|/刀p:�D}"�pYů��v�8���z���"
͘+�|�}�.�9Ė���ҶWe��e�]��e��
���+�<���_"�(���� RHnI�����LD4�0�K�*��e�P.E���SAF�ObҦ������ӡ�����􌃧���~^e2pN�P�ŵ��TyQ�d��^��pC�~��.3Q�:��Ћ�3��۩���|e�1��Nc���ϖ,Y�\�]�#�����L9�!�zz�ᣘ�j�BPN���η����$���ř��jH^`mʟ�'�rY�T��',�u^dg�R�1�/��a�5�l��J!�\ߟ�n�)�뇪�A�s�Cn5��ͤ7�ZIT�	��*�l�k�[����o�K�ɝ�b�" ����\���т����xc�^�}v���˄P²��8¯�������]O�+-�{l��k�Uy9:�-��d�^�+��u2�<@+��Q�f�M�q�/����vc��qG�뛳�K�tt�ğ��mTӂ��S��6�p*��i���Պa�p��.��6��5+�(`�8��,sk��dL�V��~�=��B���J�� �=������{�/�MU{��#����`AF���<��z�_����Ԋ5 �z���kB�f�يi�1%����T�)�������9�QZ<����;���r� ��X}Պi����(���Jx��m���5^�p� ���)�%"l�7"v��#%���̎�}��X��xwRLq�c�S��ϗv1\���qѐq�GG|+V�=պ�)	���:��S�e�f��޵/N�YQMH�=SzW c�W�8j��zD@S�]�ڷ[P�mu�^�h�/��f璾�Y!�7�A����32<�}=�Nx���gl��Bdφg��;�5�VjO��;��k?�������~پ�~��?�؜�m���V�|���<�0h�'w� r�^!� ���q�\������Xj X�@�v�i�oB�f�_��춀	��i�瓆ͦ������l�=�q�T�)$JL���q��§^�
����i�E���3?���+��ұ��o�O��(�\��w%c�:�����c�l�Cd�]jY��?}��;��gP1��:8 �;�G��)Iug�i�?����r�|!�G���0�5����>Ѡ$�X�ќ"Ywo�%ȇ'��2&�kO"�V�o�SKO5�"���a�~q���m%��	�����*M�<�S7������x�H�t��3�P��H��HS�L��W�]�)?Bl|���A<�XtK[@���(�(/4u�)jڥN�u�`�(B��k|ڽքH�tӦԤ�dk���቉P��6^5~�?x"�����e�ǐ>�u�oM�ځ�2��%Q���������w���qV S�u��'!:�(���*�0((���* �ŉIDk,��iŴ�!���[��AH�$ƞ�9���pŇ?�H�_%V�j�����$��{{�-\�iQ$k�p/nVAz*������|Q��"10�Dm�����[������p�<I3�rF��Q[w;����S"��=����hgPU���4�>/������nui	�##�yu�6S��m��������Y�_#�d�Q���ϟn����^��_j���]M=�y���G"�;�V_������cI��'x�����$$YM����p61-w�I��N����+YjE���5�4F;�6P>��B�����)�L�/�C�UV}*��ňOw��o=��Bv����wY!<�Wo	Hp8|��_����߳Mn���y�{͈wh�'M���_A�6�-BGF�H�.���ӌ�D�r�V0��h# �BHAh�@q���%{A��;(�h�Es��e��Wv�/Vˍ������0�����?0 ���OV���F*�?R(�_9�&'9 �G��$��9Ⱦc�ݰE� ِ�-H�_x��e U�lE���*Ri}VE���)Y��!qrT]�K氝��SS1����&�˧�(�Y=���������^�����#wp��ڒb��|�& ��&Û�-��q8�k��]:�\Vt�G=��Ns�e�c�/�}�p�NdI񇩣��/}����Ų,��"�D>�� QCwa���WW�>uHm_؏��7� ��O��9��NY]���cAT��V�v�u*�?��5�����X��{��0�Yg�r!��`O��ht��@���@�_G� �����~�1�].���4�3V/�ɦm?�Z;9E��v�ְ��+<>z��k~<�^@��������n����� �"<�s;�Ǘ��DP�j�5d�X0�j�z�w���Y����ք�sf�V\��.7�2{ԅ��p�'��^�:���K�j(D7��ԛ�=\�졝�i)��c�p��H��8��{������ۗϫB-��<<u��`�i��?�d�衃%h�D޶��'˫Q�o�݊��p�p���m�4���R/x^v轃��O����c~ʇo~01R�
��j�ԧV�ݰ�5U,@}۱��6��d�@�u���6�+���&CA���zw��[C�k���W x��R��?w��J咇�I��c}�d�<�1XMpK�ϧ�J����H��pg}C��U����^*WL<D�f�8��@~�1�G�^4�y�?���Iɴi/�!�1Q���r<�E�@B����́��n�O�*wte���k��u,����5���*?��.w�Gf|	Cn��K_�y��\'��z�(����xzst���u!f��|����^�d��ߜ2$�2�G��;�s~�O:g5}�#�p|�,2Jx͠"�f��81Ω��zP2���*�d0h<�o���3�O��,wsp�~��z)ăZ�tß��j%`%���ʦ�)����J�A��	����k�˽GkyFsSeS��Մ$�f(��gD'+��> �QW���W,�5�'�=S�_�ΊԓB훺C0y���M��ң�
f�5U{2`�`��6*
�Z5��q4Q^��@��ڡ~��9h��}14gZ�!z�Z�`�n tЄb�o�r�4`�uj����D�3T���� �����"nK�"��L���%;�;���|�~ڎ�͠?;א��H
�,�&�|����q�)k�ԥ�N��l��5ե��@�9M0���F�#��#�q��^�a���x8�!X7ؚ�����N�W��9����	Gh�98}�p���a��eG�Ş�h�4�������;c�ɀ�dڻ�6��������qͻ�%2|������C�v6H��]��C���s��)�H(�#�7ѱ�Q����$WX���z�J.��v� �!����b$'Ò��|��4�K�s�����ȝ�u��z�U�CY�s�f+�b>�uVׂ��9��z�)@�����e��d�p���~��wTjˑIgH�}|@�-���GI�\��~V���t��W���Gby�J�(���h��|��Zw�+�ft!�S#�Ձwr��ɰ��g2fS��!G����z�+�cP�ٝ} Kdt�����v��
q5��c�{:d�w��-=������s��&l
�
(<Fٝ[M�`,é�T;�/����<>�.��J�'I�s����zؤu�~�����w�q�!�]i�|�gȼ����%�թ��W�b:��#iR��/澰CƦ ��uBͨ�M/�;�����\h��b��X��ҖK�����%��L��� }�ks���uO���34*����ܣD��Z�%�-J��@��c&�#U� &��\����LАܦ��,��n�*�f�-l\H��M��.�峵�ř"���27*��o�N����j:��i����� uem�����:G�Y��	��i����Xߢ��	��L����j;�L8�#����@���X�i��F�Ɂ=�ˎ��8��j����xY��
��?