XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����I��rBH~����cr���0p��x�x����d��� �����Lc:ꯖ�6�����?f�_�N�	P}��� |P�6�$�3e���v+�"c�x2m�f��*���8�w�����B�D���61������5tي���`)��߈�a8��r���*
�:�x��}�&6�E~ *?�ޞ�x\��L9(J����գ_h�Wr�VM]��Nm�j�UI�{b8L�/�z[q��M"=��)���@~� cp����[ʝTP�x8�����9r��Ґ`<ή礗@3-��N�I]x��Q�_��1����[�-ϲs�%�Qd,�8���Y�g��nqSz}�����������7��!�PL�H�t�ʆ�0[L|������$��|��aYW���;��߽g��vޑ�8��>�;��z��A뢰=�.�s� �
?�]�ef\j>˺�'ثT��T���e�;� \둃�(|���KeI^_���.=�u��kQ8��%�8S�ʹ`=�0�nXF-��bmw�J{��N�#�y���1JI��`��ڭ�zH!����'Q6B[��Έ�%GT2�V�E3��6�H�+����v�U�n2���Gt:cl%�Ӽm=����1��}���~ ���F������qUW�(ܣ�$�:Òa�����Եo�L�x�kr�����;�_�r:�v��.�xH��g���}�4m����qUB�h���iM���p��`�?�j��٦H5�~�R����$�XlxVHYEB    729a    1770�>JZ��D���Ӵ{�+�TU[�}	=T3Ǥ���2�ww腎FZϼ�q\�V��3�F땊�2v������3�I�:��ע�Qm�ֿ:����9K����y\�ܒX�eܜ��.?L��<�H��<��>]����@��0*c�w��.��U{����v��H1�#��}��@�K�ڲ��KhM���|�!���V� ���Bf� f@����t���f�뇏� >����j���o�L�t�+~G��\8c(���S	>d]�:^=�3�C먮� U7��n����ڨ6�+���T<�Y3�
O��z�V��Ӯ̷�N�5m����ũ�;#��NH�+�#)�  )���YA��a���أ���<p'�Ù����U
�g�l	J¡nM8�t����C_���Ϭ��y5�I�J'��������i �ެ�"��"�����/�//��[R�r�l�PK)k6�A���	�B�%vs�	���󼋕��B-�l$g�����"y5����u,�l���
6ټGP:�*d:��Z�1�Բ�c�ɚi� �p����v}C����������n�M:Ț��9�0>zF<��D�����9iO�� �J�w�d[��N������[gR�!��YU�9�y}�.�P/7=k�j�h�cin��[�������o��]�:�rc�O�B�]�qA����3�q��ܟ��S�,�9]�l�:O?�<������Ry��Y��W����{�.Ip�'�lj1����ȉ�t�'+2�ONc��Yp����{�>��܅GW*�#%���4w���A�u����yЀ��!0�Lo�-wm-Xf�Ө���u�>%�I�a%��P�X���೽�q���Mՠ�m����Np����Z҄�s0+�1�STe�-
ų��z�Y�V틧<�9s�rbå�( ���4͂�,�*(g.��E���8�U�Ғ{,b�9�Z��8G�ϐ�D7��ƴf�m��T.<���G;�A�t=	����p��u���V�n�D��K1�V\Ư��_�E�^��8
�+�T��ۅA�E���ZN�������j����?G1Ϋ�-�̬��`yp��T=�%�sR:.�MZ&��B���X�b'���V%�}��_������)��y��I_m͊����v*m��?����62e]�~���XE��A'�_���r����+����J�6񯚺����v���X��Z[hr,��DjQ��x9��r�ULt���'`���$���2�&CXjv���.���#�4��G۶lG��Ԍ�]+8y�=G��t8<�S�b2EK,o���m�rp<���Nd�i_���+�[��~�/���q\m�6��tt8�lJ������P�]�F-3������v�J������c+�����O�1�KVp=����e��M",�"Ь.���e�1%��gw�ϸ��Q�'���d���\3[�M���c����f	z��qM�Q�z�[HRӳ�"������T{��e���a�:�:�Z��3ܨ�1�IjZ���aԛ���hD:�=��_z
,�x`_ ��ȇ�ޞ�� ;`E�,���z>{s�0D/�cQ�J:ޭ�6[c��,B~�������ҟe�a;F��7vf���R�6u��h,N��O8Pq4�E��?G������RQ�빙c�N_'�ƨ?�vu)<Au�p[á,r�2�Xʿ�Z�8rM��-Gz;����,ݧ/��pJ�[a�L�;�
}�<���`y�z�&����D���Za�P�;�9���v���R$<�:!1++9>�B�U��Q[%ݜ�9�%�[w`޼�ꗇ��#�/v�����"�Q1�!s��T�W䂛���j�r~:��ʀ��G�Z�O���R��Pm]8��,0���'n�C�A��%.a�2��/�N>{�����i~���Y��D��{��u���\=[�V\�vA9�G�;�l�k=�NO�}�6�]RO2|r8����->0��񷰚�N���g!:a��g��� ��,T�$�i
(Z�hn�д����X��"�=�F�uFq�#�,x��S�4N��J��L�O�,�n�秆�2�k�M w��}���ϭw�7�1Z�J�׬)ϣ���aTƮM�yǤ r
a�����İ/T\G}� D̏���^�B4�n��s�`��3�T�t�*#��2�������1B	�~$��j\�X�8Â��O�R�SaLuN,��7�\|Q3�i?(�L݁y������S���Leq�G���"e��)�8���B��s�����Ak�P@�6[K䐷0S:��hx[C��#��� �������/&@3xא|��"(K쑽k��x'B� ��u����V�RIz�I�=�骟ºކs�W���C����r� s�	 �q�}⮦'&+�#}C���H��?A��!�z;�_�m��f�ݳI� '�|;��ډ�;Xu�7)ט)&���Q�<[�w�F{�g��Ϛ��c��>j~}�5~͊X�l�k��Ӌp��kqg�~���Mō�ER�3�XDd���6�{�3Š6pko����o��\��T������Ѻ��c�	U�"+Ԑ��j6u$�HSB���P	�C=������Sf����6]��$JE��­�?	��~o�9��x{�>
�����}q�~,�V9��`ޜ'8�F��n{���#Y`�S	��6�q~V���</�D��"(tK�gV$����a�N��ðxĭ*~a_t�[F)��J�-���9�c���RZ�=zP��1�x^@0X哥[2���M��RP��AS�X�@��j6po��w�!�β�O��ȇѤ���� ����(�ݍ�J�雱N;k�&/��$��lƪ۩�"^���$�0�i��\���)Zu�@�`�L<��\�T��sF��r�:O7��B]?H�I�G}��	�@���%{Ӿ�$ �q�q81y;�)�ϕ����@���T��A7	����-1�Fs� �^)�]���t F���hAb�/{#���A �os���(C8ʪ�\N��Zib,٭�ٲ-OP���ӵ*'��[^�?)m�}0
+�(���|���u�zѻ�]v�S�wȗW�0d��2�MQ�zu�oY���Ph�Q��?ڈ��6��A�[��3R)26��s���d�g�CD�����YPY�ԃ\��P����6��	m	�%��Ã<+�������_���d3k��^f/:�I�+�|��2�v��ޓ�)s�8���4Rf�K�l,�*���Z* 0��D,���_Z��Wp����.����� Y�O�a?���p�"���:�>񒈞��K���z��g���+���\0�C��;��?t˴�ƭը�J[|C*#5��~����uݏ�� ��@�FwB�\y-�2/ n�R����zRe]�ib���܇ L��T�kDt9�XG�q=��R�Я*�-���*�����9���g��s8(N:�2{������P����0ɍ�|��R�+IW8���/f{��e5ACƣ���㟎�K{��}�MKʹ7�y���I� 0�v"�@3�@-\΋�t�l*�zs@��Ʉ���}�v�������̅j�&�C^_����`!R�H��@��R�(�M��[~r8�(Iq�ޫ_��'\A�_~:Tr��83!������3ޯ-�H�W�\nl�d��/?�*�����H���a���wQ]��Z�B�q��,�6iUY�v8���r1�w�Ţ�����Ϛ�d�����'�Y�z������f!��Ć? Q�R`�����J��
(�Q�3��qa��yY̚�_.e�y���vD���q�e�q����&�Ho�j\m<P H���dB��~�����?)pr��I�%����5��-�6I�b+�Ҽ�ڏL;Æ���X����AOД�,����L���#iU��ta�q��M�Nu8�@�{A�.��+�H����XI�1���j�Y��'��
��q�����9l<v�_�&���X�?}OU�i"Q�Qߨ��P�|W���C?��ǃ��\y��
YRb',h����ۊ�1 d����R�E& 16�k����S6�^��O<!�y"��F���O���<ܔ�j�yJ,�;A'��f�7��� �$�@�������m/����󉝱�ܓ-Æ(�OJ��� P�\�
���/s�b�ߚV��m�2(����}�V�S'��C� b��P)������V;;6^�ǥ���`��>%�	h�a�|�T��2��R��tf	��
D@'$I�wcZbk��?�0{�v��,�$�ܻ�P�7�2�&�\DK�s�R�3��Xbճ���^L�y��.�W#����������bE�:�T�����fMi���Q�Xv%�l֍+ϑ�o9��L���\A��"�jlmې.1'G�X%]��`L�k���̑�5�"�\"�TŚAI�����GIwy��ߥ�U�ߖ$yּq;����{P�dnC
�%�P�O'V�o�AN� z�x0��i�I����ϲ,��(�7�6�4�o���f��z��Xx( �
C�ᒇ�d)�+�1]�~��6|U��G�B�8��,�����;�|&�?!���w�R}��mz�8��T�2���~SS�ˑֹv
�HK�{��ꮁ6?���ZPh��\�He���l-�����fdg��j�9u�>}�0�� �]p�!^�p����#�#E]����a�l�ס �n�A����6�%V5�I�_���ޗ�j�#A|r�I���5�����З���}	.r� �Y�-�4=R��
�W=�:�({������a�O��& .L�檻>�&��������F��j�,xp�a���EB�b"���ptD�e~�L��X�$�R>З��`)5�u���I��1��{�����,�l��[c*��@����l$GO1�cܛ��:��ȹW��`���L�tV��U>���VpW��t���5���N���a�+�5�T��)ZZ�i\������R<�~�'�����ro!�Y���D��݆�Wl���	 �]-� �$`�]a�f	GR����3��t���.ٯ7���l�}��Ց@"g0c?��b����p��8��TlZ-0Ɍ�>�u9���W�P� 7��:�P�@�a�L��_��I���1���)r�E˫.�|�"�p��$�t�*e���A��DCE�^US���@.��rۂ�3�Op�BC�@�?w����XHdZ%�T�?1�k̩��;���R}&4��,�h�S,@����"��-�-Ϙ�+
J+�[=�S�j|k�:v�q�./�ݨ�8��*D���H�Q�.�V��y�e��Teޏ��z<����2�U kS��-�R8��K�b3�#���*PQ���?���(�,!P�+Kɟj�����
���;/`٪C���3<��N�/z����|tsX���Fՙݫ���1T����X�iy�^�3�_&�9Ld�y��Qj��l]��YObQ��@���(��2�ߞ&,��k�����?�iO!(>Y#�I�Q���|���n�1�6�~6���Q�щJa�4���8>��z�fk�_���O�n��P�r� M}�6+ƅ�P��b��]#&PBv崲D����Jr�w�-u�C%�kH;P�'9��pp\aNC����\/�++.`���D�)�.z��&��Qq�H�&6aR�b[5��)VcwдE[�j�%�)O�vl=._:��mȥ!��x�衆�*}�@ś4��w�ج������]L=��g���v
~@�%FD�×�̝Xφ�w �|H ��[�|}��^�������� ��o��]�cq�Ǻ�Y!�Uxm�D:z���=Q��m~*��S��v�G��l