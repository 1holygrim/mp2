XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd������V�k��� ��v��;�M_�2��O�K4�)n�EbP��^MO^�G� ��ݽ�v��q_u�#��ǫ>LQ)���)��>�*�s��M��N�?R�HO�c�Gg�Z�����1�\1�8���F_:E������R�X���G��K��8�pݻoGk���2U6��.v�n��P�y��4X�]��m��K�C|q�@݀ނ T�`���ѿ^ѓ���f���W#�QE����X��tf¤b�<��`�����O彾"�N6%IY��)��N��f��YN�q�0Z?;��]J��N�V϶�Yx�p=yq���/� �>z����TF,X*��QvU�d ��Ԅ
�Y	�77q]�&�b�Mqj7�x����_8��S7lk+Pϐ�VW ���T�,_�7@o�j҃svrZ�4������C��/K6�Hv>��o���$P�+0��u�����fw�����"1��TJ����C�l���)�Z1���g�K��6�ߘ�⇸�;ʈle����8D�赇[�	���v���ZW��Ʉ����g��"�FEd��	���v��.Ej7��q��M�*u���X]��%H�n�³�+��<��Z�y���M�zCZx�����т��}��IΆ����x��qo�:u��q�;�-�h�.�
J�`0�:��5�1����_�\?*��oS��F�P����+$��-�Ҥc����m�ጅ�qПdC��ǰ���t��~� ZǮ)�Z3�$�&>�XlxVHYEB    3b09     f80��\g{0e�ݭX��/Ҕ���Jc`�.
GD��Fs	3^O�$�>LZB�O' �Q��3_@��\c����M7�+�$�f�|r�v眅��}U�DC������+@+�b���$U(j{K�]���ִ8jޔ˔1&��=���k�\J�%��;��D��O[��=ޟ��
OT���.��>�}�m�;�	%J5O_�2��"��p��i��3��|��&�@���"z�X)�a�֩\��]�u��YӴ�����i��b��~��M��>$���c�;F!���H\V=����Ųd���JƒE���=7C�K�z��;}z�;����V���t�����Ϋ3H�
��j��3�_�4%SS!�8H�#�$7E��F�o*	�=��a%ដ�7d����+��j��d�CKD�+�+d�Ĺl�c���Ѱ��W��O˝�����*�Dn���9�S;^י�a�<�������j��I�Ju��2Ʃ����Fg!7n����ʗY٫B/�Uvn`����3f��(��~77[<;�G��Q�&iSw���c����
iH��A�>���to5�g ������t̐�K�1=n��l�����*�l�L�b"s��X#k��)[\�=L�CY��X����-�a���0��Dk֧��w���ی�BU��5����z��VV�a�|�5--k����y�i[��ȿ[`�qn @��β�h�M�`���wSټ�R���&�`)�;�*E-��#�[�Bn@6�w,�27�1E�EŒ�u��j�-xz�(�ꓸ���)r"r����y����P�~H�禯b8C˜`.��t]�U�.���U#���p�k����
��=�ħ�sG�C�0�ٷ���U��uJ��k��%���}/�֫y��o`]�.T˰�����j6�^�I�nLҕ0��]h寿�Z3߯���{��6jk�0�0�tS檯�Ha�1,�1	��W+�_��E�qrJ��U�>�6���X,��� h�M���,q\N���e>����F���
M>`M��~�L����H8�Z�-��g˴I�gru���ˏ}�'#�g��Ih�"23���Qb���/��.ō:��M��4C3U<[��"��J��[/jT�Z�����9��y4��r>���ʣ/mC�_�R�-��h�g�ށ=�jV}�z�#���Ml��V�F핍Vu,� �׉���J��:˦>�IY���]�I���>$��"#	��R�+ϵjA5�	~�!		ku��L����+�,����}}!�"w?�K,U���M��5D�8�Yiv��0�W��0���7]�ʤ�{��LpaE: 0���^[�W)7�O���5^���?1N���o]��d5�%;�	���eU�(n�0V^� Q#|��fK��_�xvP@#��*७F�c��T(�����x`�7��"8��a^W~G	��6���RֈƲ�|�t]*7f��PZ�!}f�e�,G�j�FV/f#�)�'�pֆ�Tu����tu�D �
�2_�.���R�~�J�Y�S�m~&�]J�Z�_0zě��i
U#�V�͎JZ�%s�K���<]Ӄ��C�e��Y�S�Zd��'�<�h���ۆX���A�m��@���ɐ�`��|M%�R� ��@��T�G �8��yH��B���S)cFkR|�����T��gA�.�\'�
?QpQh�x�T�R��QE� &���J�[���[N��w�)ש"��@|��B�q|dm7�[Ӗ�M��W���s� �g`���H�,bt]a��xu��6��G�hF�<�RUA��x�j&a����s8��Dkkj}��r4⳾Q�����v��.�&[����d�}� k��e�j�c���G#�IH�d1�)��c���_��=#dN��+f�i��ݚ=��
J�TY��A�p�@\$��MW�ÙWt�d���xf�r~�0<1P��w�\�C����[�N2�=^��-z�Y�@Z3���s�p��.D�û�;w�R�k��&,tp}�i�n+':��ͯ��{qK0�?Oܠ2 �Q351Ǽ�pWwS�/��3��B}k��?Ӏt"���F�F�^���,!)��8�# !�%	�����W�1���;
�g��m�nebVٛ[���{
�)��
����8��o]$6i�h���W20��u��w,�pA��΍��X.��hh�1� �U�-�nz,_OQ�=�!��T���?'��Vg��}L�;�)[����y�}#�;BZ�&n<�4�]�Ӓ)F���ef�rjp"Ky��W>���.J����*��
&�E�����?�JϨeF����Sp  s��S`)�¯�C9Pp�Jn�в?��gI��cK�k���0�]J;��ݻf�5<��&'Ddx�ȨP��F�H�B�����$����ƃC+�{�C1!��2Þh�E�aҕ
�������;���d��ql� �9�N�ɇ���W����Q�j� 
�c[�I�;X���H�y*��3A!�>X��+��V����`bgV:�0�Bk���r����Qs��6E��5�G�BRQ�ޠ'���g� �8��;��	U9g��/��KE��+�t�{��K�f}(hGN	��+��<T^�b��_6���e�6�t�L?�j��q!�`�;�~ȶ<M�u~n:�B6��6O���nYUu��1��5ڤvQ���j��
���E�ļ�U���*9��P������9(f�T��i�����w$7H�7�Sn�׺ ����e�����_�Ѩ��"��G��[�����(徨��5XZg�J����k8*f8�1Q�(Y�����������2�'JXOxzT��]v��qΦ��\�+�~1�e;��;���L�1�k�N�bat�O�r�����B��m�i)���'��B���o�M'�0]�'0�sW�+��{���
uFʼ����y>���	�~\�s+rm�8�s�y3,�
��F�G�4�pX@�;���p�(Sg����I�<&�K�$�|c��)�3u�@��Aki;y2�K�Y��,@�7�Ȋ�4ed�4�g�k��A4�.B�x}��}���x��Ie��r�?s�XJ��%���h�RP��^��՚��z�>�pU��)�y)��w�}��~?����г�g	��υ$���W���E^�!����KB
o��r��pnXf,>U+��Q��	�H����G"���<@��_��iG���>�E�D.J�R������$T�)�3�������T5u$�*b��:�/��&�;�/<�ɂ۰��1��nV�!5j祉c�p�*�Y��~v�R)U�� �y�����c��&�@��~�R�y]��<+7�ne�Q������O�0�i+j�u~����8�o-~�j����2��1_��[�9��!��p�`����Cu�X>�r�����y��	�a2���`�O[Y���L}q�'������(�@sK��K Yf(6�����(�`R͐�7���:�EfpMy%va�Bl;eꜛ�Ccˠ��ޱ��5OԄa1a�Ս��@I���] �HV8�0�s�b�����T���w ^���ƻ҉)X��6�-���
��r�n�[�Ө�sF�#.��˨L[7�,��䑴�����e�?���aKܩ�����s��9"j��5�̙�=���A�az�e�[%���c.�g }�6}�lU`�<�mIvk4�,�@�s��E=շ�܏M����/����+�T�bW���?�Lw���'aE/X���؊t�~Z^	�SG�C�^nC-~-g�
eש􉺴�n����E�2���y�����\���G�TlY�e�� �I���!��	�w�U��2���\k��h���"�F,�d�1E󬖩�