XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��s���o׹�	���b��ۉ�fNÿYTΗ%
�ѕͽ&|�w�������spv�ҹ
�(�-x/I��*�9�����DLɨ����agf��N$s1�l�w�x�zV�����B��س��1����K��*G�+G��Iw��"�Q7�sX��Z�n�x�=_������.���![b�"F�a�1IA~�g����eaR�
ᐾ��ŕv��1ϊ���+�(o�<<�2���1p.��J)���H��~C˃~N��^9����5Y�w&���͍[D.Dy�N7><�.�����۴+j3����(�*�|�]_ek�FQR�nCT�ji[A<�W�P��Z�ۍ7eE5
'ѲL�0\�$�uaޒ*�g�A���PD��ϝ��ĩ���X��zV8�.���VI'w	����Fo�����7̏�o�
<�PZ�UAE���(���F�����dU�*�=�T��v#n��M^OF���6���
H��e~��ꓹ�f���D�t__S���4�m�M�/�!�7�7~F]�#�<�+J~*V�f��#�b��~4�_+/욻��
t�5ޘ�#��-1ɀ��I���G�ƍ
�s����b�:4zS��ۂ<��ȷZ�Q�n��⏇����8@I�p/&0���lHԽ�Vy��������{5Q��8+����~ 1=���4��=RȌ�����"���'jg�9���e�c����>.��Y�x�+����[��½̗M�����y��u��N�!_�%	Q!��mK��XlxVHYEB    30cb     bc0H�@J�c���y�U#q��\��|�c���t�q�6i�����ԏ��O~2;��Y��:�5��:ڭ\��TL�~���(9I���W夂��yKF�8cy~�2�����*��Iq� p�Ғx-���P��`ᰪU�\��{���r��a�?n�^{e�֟�IyE�o�錃+Z���t��eӷVu,��* �跍m7Yf~�h�D�3�_��-Y.s������՚����lB�7�d`ZL��Q�6�xJ���q?h�Bsp! �Y�ha}o���^�C]�U��cJ{c���~-0XnNx]�@��Rn�[��sÆă�F�A�k%�vzNO�K�"
k��� ��%.�ǇW4�4���9�6�y����Oo�wZ��T�cn��P�@:�[]A{	q)G}�Cy �@������p�|�8��s(J�H<�8�2!�AF{�9@��w�E�#=��z?K������O ٰ09�]XhŘT�ĕ���/e�-��߆w��7�vB�ȃXu����n�E�i������'�&s�x�&�` ��qS;j^]E��#'��7��A�E�,�ײ��YX�� {.-�Q;�a�&CH�	'���A�h#yU�	�Sm�o�
���͖_2T�GvZ�[>
6���vzƂO;���>E����S8|���P*g�=5��)��a��u�l).5��G6�i����%	���W3���\�M7�Vf�S2�y��65��y�7O\�L�y�o?�F�-nhbl������a����D�����lu����̺���*ԧeE&��o�DS�@:=O�w�+�#�՚tIҬ��6�d���Lb�&��Ǘ3�"��1�g5SyW�3(N��t@��)�/u�Ƈ�������&�Z��<j�şųRy�sޱ�����W�g����}�>�mD�O}z�+�G>�R�%�P����(0�A3���>����)�������̾N*���-���!�=
S�+Ʊ�����fI0ors�n��lct��|�5�:��?y�=�iX����X0���e�)Օ}xF���a��a���c
g�w�r!
NA!%�*�Їww�H<��_�f�#9E��䛔��k���O
����f0�_R�]��'�����H[HH(߷�<�Kb^�:\����]�xZj��p����f�*Oc��h3��1	Ձw�bj�B�U��ɘ��|9�}w���[��xНe��_]r�,..��O��8���Ņx�[��[\�@�M��8z�Xr� ������	1�qhŭtN"{��6�/r��~��b�;F<,�&�x�%Q��ˎf�ؾm�*�ϝ�BF:�-��L�I��m�)a��-�����ڢ�a-?���)�x�쟑�dw2f�\ JM�t�q�gYa�ֱ#�ʘ�9����q��ç'������̝ɥ�#B>��v8��ǥ�i�d�W�!7J��F"�%��̪7��q0�'�Iz���/���~�����7$�:��,���Y�;���Ù�;�`x�;��*�ֻhu"��	�+ʍGT�i��j7O!�7���.HO�B��G�2�����+�}lH�S��(�d1��Eշ��_����Ft��[�q�ت�����bU~к&�Y6J��S���,p��n�(XR]�S�~����M�-���S �V�)@Rh�XW�Aw?���sȧk�DM��^�\�V�i�9|��X�Wu��^�A�:/�BX"M�f�Ɍ���ҿ���#��S��K:�U�A)۷�L��_>��&Ŭ�Se�+��+2l�=�<��m%��W��9�3
v8G�����
m��ֿ�aS�G�f��ڱ=��уU����/@�Z�����Cq,g�m^5WIg2ю;t���NL�@s��h�QC��	)K���6�g��ѻdM�~�*�ss���ʮ*��GT#X#����c"�-��u�@.ƈ����cu �xi�m:�u�F�7�D,���}e$��)�9�{̍�[ L�(�~�K'�E�6޲ɧ	��9�_�Yu;úA҂|��	b6韓j�a'WK�x����w W%�f� ��.!{'���A�1�bGt���OK�o�\S+�[���v�(���Yp63B�i�,�˾` ���?Z���0�tn��뛻�������9�r(T�q��D_���Ŵ�8
t���y��a �)C�#�e#�TV�J�͗ھ��+	�K"�CZ�|"��l�Jv����YM88�*ߘ걟X�&n�*o&�g1�芼L%&��M#k\�Vk�*̻}g��,�=	�x".��='LPo�b	M�l�0��C�������_�����3�z7�N�j�{�X��r~�����O����  O�#�hxl��7Onί. \�闏���/ϩ^4h�a����Bb�8Uܼ��!@�I�Hce�m����(ڻ�><��q�Hf �r�����ޛ�Qy�Z��L��`B�&In�g��j�fn5�I+��I���`^�@l*�
j�#Q2�����q.[?'��Q/0M=v�]eS�<���}��U�Nn�>�$f����cK�[����Ri,J��:0Lep�lp"���!iٍ �wW��ӫ�i�ߦ&S��f+/�Ks�cc�%��t��u�{�YQ�ң�;'�B�ާG��f�������By(ˋ�������j�����ގ�'��S��.R̟�Lcs|,��l���N�3�p����h{��%��Ls�gR�W<��8"�0QV�[]�	���k1����~����E�ݎË�t�����mn�VĮ�$%S��E>BV�{OWvI�gbᯣ��9�o�:�?�e۸I0ŋ-~��9q�ێ�����ϳ ����@����"4w��'ke��Ry7���&�#P���5i/!���1�n	9r-�2���O2��@GU�z���_kVu����֎���@�{ʙ?�����L��B��