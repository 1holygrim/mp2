XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��D���z��J!��&}o������yt���V5HC� :��#�@/e������q��C���R���B�F-�K7��䦧����4_^��H�9��~j�'Ν&yA?4n��}\<��}en������М&f�s���P�RĢBKM�U��4�<A���i�psZ1p4<��+�J�f~B)��铻�;mˍ���&�5�$κ�� �;��þY���� C�������fQWuyK,,'g���Z~:<���Akp�~��gЛ��	l�rӣ��~��Ǽ"j��R5��S��o�n�Dm�~#!�x�|^<��[3�G�΀Q6ґD��Q����9h	���Md���8z�[2����+,�`0qD����K/#�����e��!5����.�6��ƌUۉ_}�3�NŽ���`�)�~-Ĕ���vH���0"��´X��:���l���a�}Dv�����/�Q,j�
:����+\�O
��d�@�	�4�����:���-v���ӯI���2w����ڟ��>����:i��0���ʬ��Y��УL,5U�E����QR=d��l�Y�;^S��i�M��G��h��b�6<+�ik��]���A�pU.���.�J*��_��D�D
0��}C�ρ������O�nz�{�"-X�򙬘�,[�ޱ!��2�6O��S��:�	��ѪbGa�1�ՠ�{�~dX �rg���f g�7\d8��#��~z��F\L��i�XlxVHYEB    b087    2540�;&�v��o�d��F�סA��s�:��`�WB�[m(
4���x�_A�Jٖ�"�K�_�v(�dm�M�EBr(�]�t�0N&[8NC����<��0CpQo(�D�{Ч�Y���ŵYNn\=���aR��8��s���y���v;��ƒ]6	:�Y���k�"�z�- $V<���h'�j�J�;��`5��"�;S�R�I�
q�9A1!��ȃ��br�P�m7��xt��6 ��'�_���qإ:���́���@&�kFJe���J��o��<��5��z?�39޳;^X�ZͿ�&4�#�Wl�� U)���O����Pq� o_��f�y2�I���F�Z~�l�<5���7�j¼���}���G�l�]��i'��n�e�F2I�܈��Vg�4-Rys=ƍMD��������x{���(��A�e����4�S��$�%Cy Oe�H�i��ʴ�|�ŕ�=M
����V��W8�D�U|s�^��ڇ��À��`6����j�	'��'f�)�26��;�t^>�qs,
/	"ˊj�y�9�D>�v������i}s=���:��F~)��q�O���U��s\�0��:~�ɖl�6�z$��u�p�-�ɩC�M��ǖ8s�*��7RY>�n[��)�v�DV�n�p�:�r��D�fP2�-�'�Ov��K:���轁:�H���2����҃a��!5�7vDV�����#���6�����`D�e
��wR��8��']٩�ǹ�W�������aC'�jHV�z���n����[�j�-�Wq��5^��(�ɳ4 W�X�AZ ������¶Ua��:�*~ U�5�>����2��K�$a,�}k��t��:��zX
�_$O�R�SUU4��t�G��"�C:E�M4r�[�?u6� )Ƀ��T�a���/�M��JbY���ňR(�\L�G80a	,���QzC��۪�Y@���#k��0#{F&Z��f����>��7�jy�[��讟%Cv�~^m�M9l�1��Vc��$,Ќ��u�7^�ĕ��;_�v��'��+^\�;y�wƕ�n�VdCO��Nj��ﭱ���U�O?���|+�`g�6Q]��P�ܜ�/B��?h�@���q��aڦ�u��}���O��wrH���9Bl�![��s�_�:I�������[[c�5�� �"0a�~�sQ�h9U鸒��Z����EB<B��h߷�h�w�M�0	������)8�^��X������9��C2i9)�b�V��TW�'�*��U?�|�=}��!�#�4 n+�5�/S��$��PL����<��_�*��,�$P9)y��r�id�q�]E���x1���� ���9U^wZ�C���G�%"�9��u�*D)E����v��3N��P7�5ة(g�Vu��\�	�L�#,�J�XІm�����PK2j���ch�Ϣ�a�Q%
>�c�}>V�W7^,f�����~iF��(=� �=��[��<�?'Af��S:t�N��B�">9V�@����x�4�q��4� �~�3]����'�O=nG�a�9�'ekWLC4�G)䎝2���a5�V�@�">�vK�7��Г��1t�YD$�#6�����T�Y<���4`����K�5u�E�4�!XA�w#P鸞�Y�<��ਥ�)wǤ�K��V1$��!���C�]�������/�����U)_hg?��Y���`I��Eg��)ɔ/��7t�|�ҡ���f�Xy��ҭǽ��J�Tw�u31���4g�mG!K�D?l�OP%!���wJ]���#�J�jY����L|�E�u�D�w�3�۵�a��l���W�6�I�	 �8��*�f
c�8����;}f�����hh��SNav�.o�@���#J]x+j��IΧq۬���l���/�g⡶!�AzI4"� 9�����;rR�HS1�p�6�;^��895ؚ��U���3������~$�At.���������D��w�=ұ��4<N��?Ի!�/^V����/)��.��]E�Ԡ����Q�4���@��	O��/:`=��g��:G!�@���w���D���n�xA��n�'��O��2[���w<jʱ��"����2EV�t�Ր��E��ƛ����?���ҽ�`���1H�S�zp<h\'�>�~���ƪb��B���f���(��Rv�a!8�b�Y��9c�1��/翲�f��P�L�er�N᭼�&�U=����ĩ	lw����c�К�B�C�I��Uޤ����{�|�zS�P{�n/����ؒWp��˻H�����}��Q�k8��'��&e�g�WM�-�D>��4qS��&�}^JP��:���sYi�3+NHz��\�� a�疦�ǽdĊ|�{���_���C�|���Ȫkv�\j�xMN�H���Կe^���8{cr��(� �u[ӐM�������H����|pb<ΚV�f0\�����+����3���c��8>F=��0J���a���RI��pR�����[$[Ȥl|���~/�*��.�����<D^I�̹;Cܼ;3.�����G�� �ΐb$2����T�����$�kN�8!����FԖ��F�-�0��&����]�p��=�Ut��󉀐o�D��<���.��B�y���w��g��$��!�A[�tIN�Mt:�DC2ϒ%oU%T8�2~�?B	(3����l`�2�O/_|��P(`p���4�G�ck��i��r��O�a�6��g(&��,l�k������ao��僨n@E5W�������G�KCd��8v���R��-6җ�`�'v���Ah+h��̴���i~�0�i{%�D�G�|�l�Ov����7�=l+�70�Cg[4ɡ��[�߈d��%~`?�'�]#�L��"[*#�+D�EE� �W�q�t Ґ��v��3J�]�B���<U���Zj��Ny+����QK�$4�l�g�V�_>��,_~�\�b#������؝��)H=�k\�A��@q�U0U6����2�]UT�#�j��+��r{Oa�&DEfS� �Ϩ��M,��.@d�V�0z�2@ΌVN>�F)�Æ�������]��304�j^s� 	��q.C8[&E�Q��.�W�ǥ�d�)=������n�Z��`�K�g�au� �gЬXd��>uV���|�g:w{bQ�,�� 3��kW{gLP�&���B��>��P��P�x�q;�����v�(ʳ�6u�:�E��T��Mѣ��Y�\�|��1܆����&��.��Մs���%�tiYZ�h1���y�&D�:Tuy.���X��!�ng��@eƽ�@i.�1�9�V<�B�˷��\)�>\�����X�W���F����/k&���}��Ku�0h��9�����Y��M���\6�hP��<=kbT�.�_M�٨�����-�rdS�+Z�C�(�P�ud#M&�P��l.��9!���`s�"�m���
7�	<s{cb�r���<t�̈́@��\����ъ�bi������$$��s�2����­ߴ�tJ>�h�/	��%�ЦAP��/1�*ct�	���P嫮�V-O
��]�Ĥ��%i~/�W��S�k�ۡy�63Qw]r#i�:���1���X�����B*t%&\CX@��YB��UDA��CS�ua?A������9&�A�M���\	���\z0�iJ5�t�&Pelw$I�$Qa�0����X��f��5s|�ϯ*�6O�������;�&j�R�R��i��Ov�Vq"���>ct�K&��#k)�R��u�� xn���X�o�qU}��	���7�� ��dj�t'˂�:���v��gG�ޢ���벸`>�N�����o!浤�{�Un��bX����k����*���[P��Ŗ��g���m����ZO�G�@3?�]���5)O�Y�F�.f ���������Aa����A���lT�>�H	�pN&��3Y&=����p��"Dedu��BU�"F׾��fH��uKzw�4��.	\DUG�u��E�oК��	%�"~� ��rf��f׆�ɗuS��S�#����z��_��YUa���pg�7t3f�GW0��/��dtԖ��.ՈS��B+I��5Ќ0{ۣ���1O|���Q�cx0��
0n��=4���[(�t���w�9�85""�f���M�_u�a����m񬀨��|Y�
����@#����#�n3����x�tR�*�Ax`M�ɠ\k{-��|�Y%�v-S���\��T1:J�ߵ>��Κ�'u�Zd��("͢@L9�6�2���e��"l�ѧ�����>o��B�� D����t�0+�Bx֩:�ʹ$��mO� ":�
�z�)�ܟ��qNܩT�;s�^e\����(1]�!�a8���x|�Ƚ���[O���ԝ?��4��#�ZR4
w���@�흠wM��`�"�,PVڦ��@Glh�G� ޥ� �[�8�}�?��z�Ԝ<��(�Q���s�j=&a;1��TH���er�NJP����0�������:��u�A�}Q�#hL�4B�U���ˊ]����P�#��Ȟq3�ƗC'�x���E�����M�3h�3���H*�)��-��sx�Xb=pN��(-��An��'�7l���bJ�����K"B��u֯�n2�((	��p��'���qo_.��'�{1�1��1։�x�9S�6�{��T@,l��y@P�<He�E��t|f������)�Mق'a�7؋!(��߰k�����Qׇ���6�����苿e�����@�<C�4�`���%S��e��7)Mƪ��Y�O�6�yUX�GG ?/u�3WN<��U�C݌ԉ"d�^	��;���*���%��p�~�KB��g���(L��xf0a7��ZL*�.A������D�q���x��̤&Yd-�:9��E|pˏ�nc���c��?�s&�.}�0�� �4����k]Y}�l&�Uz?��θ5X��j����gg�B��1;6��ro� 妡$��n~ލ�Z��fi'({�w�JOPM4d��"�ŕ��mKRvb����Gxi�����B?���s�%�.y��?�������Ԍw�= |��t�wQ9(hci;_��\;��e���l"����}��I}��Jd�qX@�aþɺ�2��e� AS�t��O�,�٣�e�����a/���(�W���K �S�9Y=;���IeFC�4���ֆ�0�ÓFB�?:�Pot7�s�g/����;W���/��jN����Z�.�ze�8BV8~�p�ܭ�����
��ڑ��~\"�5rT9yMj��x�;���CwG�,q�b��Ä7e�H����؆���EO��g,d�|>�2�~$!jw�����	Z4�F�ؤC�Rc���U͡p�h�n�7�3���+F�����{HiO3�ms�����_̛����������T���W��:����:��X=2�x�N��=�T�W���+8A!��ȫ��������f ^��+V:�l��G��{��b��$�x��f���1"�pe���ȱQPNYϊ���fU��&b�dC:������C(X��~�}�k�"�-@k�r�t�mʮcN����٠ad�*& �����?@9F�QP'�5���p���c����շ �	r�#V�6E���	Ԡ!4E���}�����f���E��t��6�����K`d�b+�?m�
m�!�=|O�Y�ΉpɁ�����'}jK�����A�m;�B�{���a���L�^�['9�b>�� D��U�����$�
�6O)�]#Y�ZG��o�;'EF꜔f��O�JȻ��8�^�T3�ˆ:>٩��D�PS���J���,i���q�1�,���,�X��#$�����L ���o�>]&�P2�b��U�Y�f�n��������6��Ȧ�^:��M(�;��k�tr�(:�[���>`y�	�+�(T����dx��˸|rX�����Ǯ�xz��/C����$���g`z~��͜�@?"f���&`y!�*i&����0�gg�����9��	��d$@~�Q�p�_���t�)�9H��|�nL��D�SG��7'a�P��]�S�O����_^��\��V؀iS{0�S���Q�AyRW�YfD�֘8%��/ ez@Hl���M��l��%�<����������=>���]O��:d���Q!~ϓ�pPq2J�fc��tV�����I�i_2�Cl�`���}�V�+=�d0�T���R���uQeD-@�^����k��|�"g%��e:��SV��\EtI5����̝J]��mW[��f )j�ʡ b��&%�=3�f�@T{Q:���I*u�}.2��A&.|g~��7R}����̮D� 5�]�D�&X��!��"E��j��z�"��Q5B�NK���^pB����-��+HqV�Y�u���{����5f���_͑�9�_K`|/,g?#غ��؞��P��₏-��N��Z���(�PV�cK�^�֦����~C4sد�Z'��/-k��7��˸����2��XI3��O�M��B�K�*��<����B�h�#�:��"��X�ry�D1ͧ�l���m?���ͭ��d,�(��"���s��#�AV�X�֣���}0=�du%�ܬ�q��g���1�È�=�QI��kN��օ�n����ʊ�OJ}�qn��N��({���-Mة�ߛ�����e6�!�r��Y�����7S����z���Pg�����#�`l궿T��O&`���ߌ�c紁���?�?�������HԳ�g�D׋*�ݳe>,�t��OH&�|S-bY���f�`��U!�>F�����/-=�����K�guI ��|�X�����2т��4�H#��y��w��w���;a;!��v��Z�߱w�NrM*��C��I�	��ޟ�'{�A�>[�HI��4j�m��K�g�Z�]���h�5�#G[Z�WL�2�Q�}(�J�k`�^9o̊��8;C̅}���k�H,k���t� �N�CY
._����f�>S���ڿ�0TWO��|��3�<���^�����8�В!-�O���A���|��Wv�4��=@0�� ���)��C77�}�E=L�<EU���z����S^
�l��?��B=�V�[�l�d�
�
ӥ%�A�=<�mŸ�=4���R��T(W���kt���%�m��x�3q�Wԡ�mR��!�T���h
x��Ќ$�9�=��Zݪ�Y��X!����lO�B/ݡ�h���ڵ��|�w�`w�hۿ�(�D2����W\���UV�XԽ���HA��5W4O�j�;a�����9�%���otDOje�hk����mե;F�4�^=���m+��f�J�B|�:�H��ɮ�8
=b��Z�mIDiKB�w�bܩ|�]>�z�R�����#��"f����kD���1���'�%��/(�4"���'�sfR_'r�(��Cef��bÚǉ��Zp����	��FL�z�	<Jh&��T9oV�O���G�]��Y�+L:���!�*��i��UeLA}g�Bd`}e�X�䢇#ߝ2Q2��FQ E]�@CG[�{��������s��ПK���n��>��:���)�1��]�aAF6�[\eA�Z����&�I���{d�<q����=��X�'�-��@��A0�A\�ʑS��Z
Ա![``��sڻ<�pQ�X8gUS�"�/��ޠ��7���X$f�vh���gZ��Z�;Yd݂$�[�� B`C�$#��y'��0�Ҫ�`����Y��qt�dmVG��z�!uiyy��Qx���n��"5����q�U0�� ���e��g�G�\*��@%�*ˁ��a�m��4!'�&���m;CK���KR��pm�8��=�!77�R>(e$�6"NN��7t�{��m���}���Khp�-zX�bwU3.�� �����"��>�+��`{J3�+x��ȥ��j����B�R{G���=���|����m޴�N�_��h� E;D�<�C��u�?���Ku>�ma�U�7O2��Y2-��hIH�\?B<WNCT�����PdVc��
*�p�Uȟ�B=�bA5<���k�޲v��W\R��cHIia�P�}{M'��U
!#gE�f�4�l�������oz� ��ɏ�Dط��]�)�	9"���d���a�[�}I������hJ�@�m�'�TQ��aMS/�|�@�m=�"!\�A�oeJ��}�u��VbH�����P?(�d�e�p�~�aZ�Pp���ąbGU�L~�О@�SY�j�v#��BJ�oـ�m�t�Jͭ�����T�è��[A7�$��:��`���X����S�H!a6��,4#o�4=	%��j%�2�( ��wp�&'!�-�!M6j�P�{��!&Y��I���{��e*��G�h�1���<C�@�̴A���;��C�7w�K4d�Y�,���z�1&$Ae��>F��u��Y������x]�����Z�����Yb�ֆ�?/�XÑ#y�,| ��J���J""WsgC�pBf�(����DAq���|C�:c�e�e
@�@:�#!!'n:���Y�9#�)��޻�F}���u�)���Θ����IU0������Ֆ=�]��"2K�6ŧh�����i�D��{��%]�-8w| ��R�K@>������I�ݚ�j����M+�<�ȸ��[���W���r�MQ���k���)w2�Fp#�
j3]$����h�}��Y���惷����{���co��i���_x?�c�qLp$��P���ܚ��-5�*K*8�1W9P�i���(��dDkW񚉽�rVC�"��W�:��^�x��̨jd���kh�jmS�d=6멄��iP��xi�K_�g��]A͡�\���;�"���}י�)�_J��1#���v�?SFک*��/���S�vj��6�P"�Q�Ǣ����3�����r���A��7]Ur�O��lTӏ��LM�c?NgQ��6�O{��<"�݂a�Yn^ޟ���|.y!��&�1C��v���K%���N�B_@X�G�U�шAn8/yZ��^ԝG[�;Yg7�`O��d��P�
��R�d�hUJ�KC����mbRi��p|pL��Ch���t�%J�g]֦���{:������$~�)	u�ڴ�f"���?�Y]Gq�mU'�E2%��ҁ�'A��1<0�+�UV��"f2衃�T����`|��M%w�}}I;�c��cQ�ܮ��\�����%�Q1�a�U�ts��CG]���s~���-��?�WZE �P�8^���"���0�����������sS��