XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����}������Ҁ�H���A�+v�`��f�/"����bt��+[�a�l��ј�(�QPy����,֥H��˘[X��8J���v����/�x�K�q;#M����=�!��^�A�G����
�_k�{�s�jݘ��4���5����Gw�Q= (S%q�eg:�Mώ_� ^��p�o\&��ǂH&~�q�?b7�8��_�uCv�|T:d�]Gs�3���zl��ڞ��f��Q����:��ʪ�;j麌�KF�OA�M~_��f;kQ���儦����"Z�Fbm��a�����J�ku�v��Ǒ:��}���R�ӬO(�bIɈ/�Q/�� ٦�R���/�� HeZ�LyN5��Ͷm:Z�W�nGԫ����vx񫗌&oAڮ���ք�9m�
I;�{3���s�B�N����eI���`$�Е���d�S�����X���Ac;��Ƶ�رoX��/�3=�m�gZfkM�5ǫL���0AO�(�2{�l�"�asg�Q�q�� ,�L��F&�?��#�0g];�L)��D>�+*�&L�����V�
�p�� qJ��셓��]*W��K�S�����<`�Y7��խ�$��E�(�gi�;Y,�Z�n�%9����ى�\a˶���6���wϼ	���xJ֋)������Q��FS>:�|�JlB�V���/��%)�M��X����:f�)i� h�Gm =K�D?��g*��e�	N��,�ʋ��d�o�dH���&XlxVHYEB     e07     680�:`=�$�tӟ >}�6�
��T7I/��.���4���~��R*��r�o���!�aD�����YHX�q�e40���E�f	)�%es�Z!�z�������a�Tj�Str��b���<��T�.�h��G��p��i"�p������0��<��*�}����ׅ�7�L�/�꠩�ӥ^MaK@�
k�m6t�f��Cj�O+�I=��iv~�!�/|J�])�d�g_�_�J%<����H�C�q�r~��mgğ�~�h�����ǟ^�����]�~t�*��[�����2����r4�8�v�?��F1+��uMF�yf4�#՝$��=5����^!�����Ύ�O{O}ߺ�����.�H<jvA�	�G���Q���q�� �nY���1�5я���B�k��;T��KkP#�L����T.�úUd\-5w�g$b���<��s���9֫'2R���כ�jTl��}_j���8XP�##�#>)�"��K����@��vT� L-.�������̓�Y�-V|d�>@�ǠCX� ���t����nѰ!ꡓ�!�T���d��xw�ϧ\��P��a��Si|���Paa��ȯ7f}���øܳ'WW�)�aAj
�,���5G�
��N��?\�Mv��bF3`���W��1����b�Ӆ�Q��}И��Y�J�t�s�Z�X��r�rjOe��#v�˓��y���O?D����!-R�����^x9���?��K	���3�%�p��azHP(�>[N�+괙)�l�F�p�;�gO�
M�,��(�3<`<NW��e�L��r�*������P���]8^KWF����Ѹ"��OL�yGH���q�
)��ξ��:j9$TF������ ƕ#S�-#��	���e��������u?Z,�H���1E�rs�4G��d��$��P��v������5��j�!JΛvl�	�����
��\-؞]�XGn�9q��5��я�x�& �Z=��
x�ON�U�BV���L��s�}����O3�Oi���贝���zV�s�ti�SU�v�3���s� (V1�W��ӴU{���8� �~5��Y ��wY��$�C����T�}���J��9Ӳ��4�sW�&;�����Gt���CV��D������F�Mؕ��x�a-�e���td�&R7+^կ�3큉�9URXCK]d�#-o1V�%au��Zwb�R�j�9���H��^�<���ƌ�lU�f(�wùE��V�s�!V:�]͓},s1Gg��ݫ�����ܴ��O4{j ��M2uπ�N__��o�4!�OF��j��c���+���8�ǒ8�w��&��߰d��JV��m{��W��nT���?���k^��L�C�xm��t!���S'��SK\")N�����@ ��;V�m`��^�Ƈ<!��x���hF`��K܂��s2���4�[���N�bf�d��1Ϟ{�u�>,��uQ�F �p�/�!U�n�!T^�׾��ɳL,��!HlB�K���K3�XQ�AO�"@�FA�!5�w�͈�Bn��#��_���E�p��k�tC�V�{�+ܣ{77��K����/���R2�@���t	�i!��<�z����;*�H���t�o1�#�Q�����")@[