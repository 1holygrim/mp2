XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���p؁�Ύi�� ~l`Mt
��8=ݝa�f1p��y%�oP�#���8_x��k�W0x�?��?ƱD�������u$��ߴ�wȴ헋V��-c_b�)�c�T���{�@�1��{�09u%Хi��3�;QZ
��F�s�	���_B���:ӳ�(���74?N{�l�����V�	!�v�{����~SחU�G����8�K,����<���{���<�2�F<�^OGg���a�P��@<��.*[V��o��	��> �����z���*Ѱ�'�^����Rϔ�=+#�[�a���T��V��c��C��h2Os�j�-)M���N��,2�U���X�=�!jK-�o��4��_Z�muP=���}̨2$��NCԑ>f҉�$/fb4pQ�?x�P���1�x�\�^?2*N=����'3�+���|��:H`ٲ�nٯ��rɇ��rԖ��H-M?1zjru�v�Κ��nm=2�X�ҁ�I�fXi�V�U�0=>1��+Yߡ���dE��hA?cdv�1HU�����n¥�!m'�z�'B@N��Z�V\#f��lɷ���日lX&��WE��w�|�I>�A�Ǽ�1�I��2��9�TGNY�|W܆��TxIԔ��j�H���:V���?t&.���� �E���Ąso�:ͪL|����<���[�l���c��$Zd�0g�/Jc VY&B툟����Z���2�%KiJ�
Jzq�'_ͭ����{�p`��Tk��N�r���XlxVHYEB    fa00    1dc0��l1���l�e�}JȦ��@8�9�_C�rtʾ��_�˘�d<P����t'����V�"��f��J�u���z
�̩uR��5�|�{����,�R�ƜSS����pA�Q��ʱ�oR�����t zH����E�Q����út�5�@��%0o�}0+�7�᫋	���@�!"A����F˯�BwC0�V_.9%˄�UgF���7Y4���>�޻��Y8|����ՀNEu��E���+���ѹ�f<���X^�g��[��f�\0������ȗ�����2Ԩ�>v<��׭�:�.Q��o*�?���'��X{�abv��ǐf�KH�(+����%��q~�1`��J�xB�>�ٵ��u�@_�ݸ=~p���ȧ�aL����C����O��I�ؐg�A��##�f�ţt�^dfڕ跬������z����,"jK)��χ�����j�<�"ʚ�i��zn�	e*�V��T��(A�[I���2��E�-rҽ�Vw������(�\����%���h�ă�츫N��DR�(��u�ܹÂ��j����0xΔ�=�o���rmb��z��L�� �s>�ɸ�hSԅ���П6�F����Q��'�0/�z���5xà����og~��dA��o�9�|ȆGV8�b����I�8��ą�7�����S
h�ZP;��:V/�Ca�O
.��.C�I��b4�f7M@����]�1<�Г�0��&�m������dF=6�p~dK�>5�B���q�hm��)/Jυn�
��x.�]}2��1�����v�V�%\��sC8������)2���'l�+Hc��M����p	9��"�ͷ2�AC.���v���,�
�C�!R�t�j&��a��bL|8hXR}���y�|v��z4���*)��c���;:���(%���
��:;����F��`�LCF��b�5�����E�B�L���1�5�5�$����=b�k�$,9�R� ��7-�RVc%U*��x=n��\��K2���6U#�]�>�KaI�n��}v�"p��tḷq��xS�(FNQ�w5���i�9����x :��/H:Yb� � ����d�S-B��t�gX��t�Q�J0PNU�ۚ���;�;:��qv���Ih�<�zq��ޔQi�$�v:�;�R ����F��Q�r���m���1�㯽lTMA���^o�K+ Hv\�x4�ƷF߅8��Ġ�K�nW���#��?��=��v������n��y1sZMkSK�9XV��}΄n�CU0�ґ_����V�+BQ�RT�w;˒�#,J��F!?]K��3gs�UЕg�X�?a����>$F�J��4p�;T ��j��I��1���6�����bq׊λ~��ɀ�90��X�r�6y�i��G�N��e��ꠁ��^ҟ�`�
�#S�ړ���j}�|���u��Q�2��δ}��	����ggD��h&���B*���i�&έD(ӆ`Ӌ�]4��S�q�Q?�k�fP��䪣�Z7�`�)�g3����R�ֽ"�;]ڷdI�S^����N�JJwY2�@���P�����?G#�P,	�|+mlv��'�����@� ��~U+PjP�*���4�g7TKz�K�U]��N<k�����le���)��Jх&Qg�#�Q/hb��E%��<K����Kڨ�>���у��#����Nވ z��a�0W�R趯ۻ����G��b�®���C�SNx��ɜ�.�{s�LCG����0,67�"" �*�o����c-ٓ�!x^�H����H����x�2:d]G��)�a�:��_�YmcR{�� �Q\Y��<�ǔ|n��.C�eT��-���E*�xpŸ\4�}�z���&|�����/�����7��f�����X�.b7��B_�MA��.���#F�TV��CW��;��P��eB9{igݺs�7{���� �������Y<n���O��{UjB�pZ4J������::,��J�ț�%�a��<�<�e�{��T�a��~��Ƙ��뢌��pho�D;��(1��w���b�^
������b*��;F~��(1�L�Ѹ@V�?��C�.4�����Ŭl��R�t2ߝqCtn1��ED�9��Ү /g-�ǽ�j0]�B\2>݉��O�x
E� Li�)UG��q����*B �ױ�K���Kb�ط�Pe�*�TOy�媬���Gg!16P��
���(س]�4���i�l�t�1����k����
��U�aҏﱙq��7�n�~I"�q�%l�,�i�m��v��jX���2��G>����N�6����5�*L*�*wL���e���_��F)h�/���\��ڢ��<dܟ��lI�]�j�m�~�|�x�� 	ub��%׼ ~a�[���P����XH1���BW�״�E��Y�;�T�	��i��K.^�t��>�s<��V��
�y�R��
[�`�j5��h -Be��*�i��pi�lZ#4`kyS��#�V8l�I怘�j#\�R����u�D�gէ�k��5ռ�F��q�'��`� m�9���1��B�*d4gC� !�zwS�k�%����a
S��!�:�4��Кw`K�\�T{�u^�{���<��Rҷ�İ�ҿ�(ގYH~���E�M��HP̓:{�ۥ�;�?
��_>ŋ�I ^�E/���w�w�0��|�)��l�����m >-��/��+6�g����P֚,�>)�A���<>1�J�C��NT��Ո��j,�P2�� ha���6��R�<Z�5��SB�na�Q�����K�/Q�A���߼�/��ze��T�]��>�Ʒ�Z�v��a'Tpyg4�� ����K N�Ò`�K&ZZs���N���Xug?�������2�̄���Fh���N�`��'-,�~��J-��=} ����#�4?��.�Wh}b���T���R�(1,�mtUn��R{	�w���Gرw��~~ʽP��!��������p˒�}�/h)Y�Ҋ�!���pi��CW� ���7P�9N�W8��1��$B@F�ՠ��!�B�J���O����O��qF�$�3k�e���i9�hVSV�Osݕ��8�o���J�;��XF]�s���c��Kr�w(��:�e�&
��B�}��9ms!b��o���㳈������m������=�Z1���������CU�g��<at����m/d����oY�o�o"����'���O3�1��n��aǿ�h�X�����ҹN}�M�r��m�i�~�!�����"�
��pQ�a܇Sݔ��
� 7h7���#�m�|9��W�.�?��.�s����e������R� O�-��/�X�h��V��d��t�W'O͸���QҧݦT�=�t�6܏VB�l;���7Xhh��8d&��v�g;�+�g��m�S�*@���g��s��\]�~^�����O�R�y�S���x�QP� �3ҭ��Lx
�9�I/����<�q�A��z/zT����Sۭ�m���DQ�����'�,�_���<�'�c�(���~
	���b"�����#˂ta�>��6,���#�~�jk�	���)W�7B�#R�Y�Ѫc�U�)��s�4"�W��VuTF��|
�l�w㥃���^Kx��(��i#�}� ��;�K�<h�s��m����^�Gw����A�~%���hQ�ե���%
�T:�ؚtR�-�1�&ȋ����wϩ�Z{q�d���kb.�� ��#���:F���XJ��#���lY5 �U���Xo�Gtϱ��{9<���BˌO�;/�;|�|ၶ�����9�W�{��[�wV�.����w��e`O�V#�-��� ����-_f1I�x6��kJ�/[�6�0�X�~�TX��\�X��e�����LWb���u��P����Rvo7��l�9�NU5U�3�2Z��9R��P�!Ă�0l`y�c3T���3�Q�b��"�	�������K�l
hTip4�h�r���n+���4����ɒU !hD�
w��|/x����N;��_�jUAm�y	�]
S���jW�|>���SY��&c��N�������b�<>E7��� �ٮ(�=ݵ
^�WX6
��9P�H0l��GVKo�;%�Q\+C��s�_?{U_�Db��[��m�#؇F������亁(]^�,WU��xu$!�͑=�x�n,��?�}���C�9*;�����Js�Zz!J�Ӊmt�nw?��i�һ�l�=�.*�L�CF�&[$�-��	m;U_���0�YP���
ݼX�s�����/C�A�p*(|��S)[z���4�a`CE��:^2���2����_�o^�kO,׫���m���S`���{��\3���n��g���2K�s]`\Ӣ��TS���Y�H�z�x0p�-�_aFHy��{0��i�IK�g�D:I9��/<H��_("�n��Du�@�U�#way������ '&�8��k��S����1M��oH0�à8g�ל楥��dA�t�O1�P�$���AM'k�,}T0(@�rw6_w�������[4|h�R�`C�,�M�(��LH���J��~��,䏍m~���i)(�1hm��6������&�����ő�VRt+a��iR�Y"����AA��'�-���h9�>P2��ۓK�[|�^B�𦕤����e�տy�K�f�a�V ,�Ȓ�-l����R^�f�pu��C���
���7�����K��D� �T(\����Y}�3�Jt�(Mm�(R6Ȓ�*��dR����;��J%Pq�i��XI��w�m2G���aT�59��b�-&p=Ve��Q�XA��=���6�i�0WLVL��������'��ԫ�Q!}�m��'�y"N0�Y�|DI_Qt�i�Q��{�9��Y���	0&�SSɀ�o������������}��[��-B��iO���x�y��O�l��$x���ٶ|�Lõ�id�zGw�;�� @�j���
𜍫��Jndu��m+	1~S<+h������Yc���\�Ȑt��z��W��)�k��\�"��o�OҰ~����8y����&X�vD�WS|x�D��Yz�A�����a3�:��I ��29e��# |%7�$���J�j�
�=��7�RF�)3�8շ)�iZ{�iN$��=Ä�x̂׍��^.N�96�7<U�23�\��
Ep�s\=�v�{���hy�Y�!�S�n�
�Y���$����1}ؑ��H{wr��	A������Ƣ��#��-w܂��b󂙀�t�����'�j��y�k*f0�2�!3�(E�N�l���4��[��5Hg�k����h�F�(���|����(*K��Nݧ-�����+�g�H<�u���g|c9Jľ����$�3��r�:�ַ�/��pT���,���:��,niD����O��X���X�f�{�e�A+բ�H;a����Ā��\o�ub�2����l���1��d?v�vP�<�Prl�kM*خ}�k/f߳@���>�0���A���S��Q�����ʺ��#�%*i�H
������"���P]���?�mF۴�?��ir��`5V��!�vW��[B�6�x_S��.U�n��E�Ō7�YCS4��┹Ȳh{n������A�K��Zfv���A�O5l�Q��0j$Y�v����O_>Ӆ%j�L������)>�v�(��$�$�v��mA���/v(0�_��R�L��\�6����B�[�����&���F�b��-��7pM&nd��|�>���"��}��<���K�I��efQ�������z�:&�4d��5��1�Uͦ����8��q+�ُ���+����EkźĬ�XU�ʉ�~��4���o+y`�s�8����h_5}t?-�ge�1�,D���u�-U@K���Da�e�.4��[^+�*=��k���o� �!g����^�>�3T�b�wA�6�`cG����WGGc3�ycp0~��l�r�@'c}!���D��)�<$��D׍��&�^�v6���}w"�U�px�c��P�E;H��_�xi���闯�����o�v����v6x�H�~,�dl85Г�� �J��_��Q����2'"h��|ģTP_�x�*R����Y��
�2 ��*�g��L'ɩMA���E�����X�6�I�����=��:��� 5�m�Bخ�zp��i�q��|4����� �KOY�iO,������F�ܺ ��¢��km�4�6��]��I)%��U��n��!8�n)U1�i&'"�|��O�N�w$��s���v�{0����S�2���ϗ$?K�OS��1�#�eS�0�ؘ���S �?��鴀8ok����r+����j���4e�IJ�MT+������=���
Z\�F�CMѧ������hqS�����ܠ��>���'C��뗅������#����d͡9���`j;Ѷ��3-�f�<�2P��D"��Dy���ݧ#�%еm��j�����l!�.��M� 8�C��&�2��Mx� ����mk�#O�^�ǧɝ�@6�����)FC�)��N'�|1{P؀�Z�ߚ�� ._Kx!�)�l�%Y����H��PȴR�7`�h�UA�Q�r��Ĕ8gvOs	W=��F}����st���u, liC�z��^�<m��ޱ����Q�vq�9���li86S��z!O�=-�ov��65�Bx��������8�m/��l�zgI� ��U�z�x�	l��.�Ĺ�;� ����g(�XIMő��L.���9D���d t�4D�w"t!#
8 .���tq#H..��ֹ�z��6L�����y�C;[-K�9��b���-��gH��y؇ I*�%�F[u3�E�۰6���|<(��|;.P�����u�r�S/������~'H���
�Tq��}����ش�D �Lm�-���Ν�(�2*,����_ɝȄ�S���A����j��Rc��fê�$}��
�n�8HY�l�9�����Pu���_�4��L)�6'CG3���`�P&'�2��ORf��Ϩ3/�ff�7|���*��@B���R��=����YP	�	�~��^_�N���aZ��OG�g}@���i���K� Z�?�_k�G<�,\���� ��1p���4�'��zQB�����-�8oc�����P�e��`
}�Onż���q�Χo����p����|;
3�n�=:Zp4EfL �_���hLT+K��*_袽�,%�Z>*�Ԛ����'����������o��~��Ar�jA�L�TTx���vw�{�m'��h�O'4���b{m�Sku�����L�@dQ��u	��	E�E�Z��n8�)eB�j����;-jL��y���,\'Ii��nd�
�����M=��BY�Y���)!�x5~%���L�J��4s!����%�&XlxVHYEB    e7be     d80�}�Y�݊�.�A>M'�FZ�<��i��	o2����7J���s����*y`}*��I��5@4'���ݜ:���i4��Y:��ҾP�6�NI���g�ϡ��G���/�5_��Z8��,��^W礠e��(h�.�T����L�ݐ��-���Ɛ�/��,�&�M|ryW(N��d?�؃?xSw��e���7���iD��S:\��	N,��C"&�̜5��pZDQ�Ϸ\�-�� ��d<��3�Q1i�n��HܒE���RA�ns�;�!l+�Ql�l�uu���b�;([�_?�υ4��3Zv0j����m��d%C�_�M�ktM3b1?xK4-뭞3�J7��	�1M��!�\�=��:c�t,�3܉����R�o���Y;l�v�S$z��[x�2�q������܏A9�sܸ�%)8�N"c@� �rL]ӭ�t�J
�6L��;^�M��d�u���O��N�my�s76:R��X�����>�C�X�V.EJ�tL��и��s ~�IT���cZ�Q`u]����RUKL��Hߋ�n���t	.
{���,®1�ޯ��u�D��Jˊ�*Ǡ��x����~�Wg?у-\q��,T*C
�7?I���M({�^n�����p@eb*���OP��Pčv׽#�_]n5��g�/+E�&;QL"=�7W���2rZ�lu�m��N���h=�[�^@�Y��(���L�#߱�˽m�!Z�ɭ��4�����N����H#^�*<r�Х����s玅$'��ZW|YYj�H�'���kh#�%"�J�|B�QQwə�E����z��uK�֮;j=���!�,��^�X5�K��F���T���_j�V��7���̯u]�q�h\�v�y��D+(�z�wܬ'�!����6
�C�R��!q>���8�����\DM��"8D/���z��������g�_���
̏\M%2Xn����)}�5���F������^w��GbA"�+�p�u�o�w�"dDۓ�X|
�UM(�`|��/N8C���"��WO��f��z��1#iMĖN�S�|ێ˒P͓�F�(w������/��85!�
R"�`�-��Y:��YQA��mS�� ���E	���c���"U�~ʉ��F�4Cw��5�r����9G�-�@ &�!W9�c�G�\�߀���,>&��j7�ӧ&�Hkv ����d���� ��q���`�~!��M@RH*�*ޤK�
�5M�D9�����[O0c�1�n�4]l�GF=�^N
�Џ�}��Zd���<xΥ�/R��XݰM�>���rp��S�΍l"�<L�#xh�-�a LTm'Fkj�uQ�[5|���#�>8]�@"|%��l�Qg��I}�Æ�~�{��'� ��+C�n}��F-iK7��� pdGa}c�m�XQ�3��V6���,�rG?�ٶ�7J���D�X����(�|2� �͙>ɔ�ך�B�/�!����aѭf�)�I'�6�upeq�Ûd�;�8CXr� �,�u�������`�=/c! X�j�+�6�g�[d���a�0��˕6��c#ɐ�3�{�ծ��u�QF����qY{�&�fZ�Ҵ�-YgLÔ�@���OA���.L��9��t*ӊ�,&<�z��z����?.
���Nq��Q���w`S�1�[�cp�0L�e׆�vǆ���!.��퍎C������=x̠�6G�]QJZwg<�Ч۩���Ti'^��i�~a�]OΤd
9�f���7�����	!6�
"浼Ҭ���/�_�r��{���t�����l�p#�LO�G9t�z;�lC%�tZZi����xx��}D�n�]���d�u?�91����ߐ�����?)]�2P��)�H��
�ߕ���^��*7��ݮd,������"�Ӈ��'h�?�:V�N�P
����~���Y��󺌽��[��r݇��#y��4�"��syfZ���)kT�X����N�7+]O��΍O�i#� b���,L�����i�H�"m����˱|�����óB���d��w��GG� 7>a������Ko���0,�+���H6~8�����(o��<5կC��rix��ŝ���\RnN���ü�:��/϶��\���jdJ�X�(���Hp�q?��mO�VQExMF�S�:�x���|8����qt�-L �� H}�H<q�Gm��X7
�ؾ6�3i(���b:��g�*�-P,V?PEmIMb���,9Ρݟ�|FM6Y�	��҉HV�`�?�5�e�Z��qu(
�j�A�cv�~V�9nt��f�k�AVe��3�?�ʮϮ~B[�����J�� �=\nA�i�>+U}/�ȉ�`��wO\�#���[�?�dP#FS�_��~��|z������>Cq��+�++7��2�0u6
KՌh�f%Z���}�@o�	��2G��ӦAe�)V~.,6o�N�{����ꋺEZ'G�E~�*���sP10��[��\�{v*�G"�!���~N�<�Ǝ�_�4C���?s��8Q�;�=���;|�ZA����}�?t��T�魕�lI����@�!_w���%�O�fv��E�
��`�O8�T��m��uB�B$@\ ����"��֨O�}r��5�v}k���i�m�j��M#tr��"��������<Mï|�4x�a�Bp�	cb��Y�q7ߝ'�v/���&y��75�-Hx���Ot<�4�Y��j%�s�%�G�,9��F4�kv07N�fg�!�cn:7;W�-�/�gJ
��v�lf�Κsҩ��ީH<�+)��
��^N{|��N����/�c�o�<��)L���6�3ֶDx�Jn2�"�m�gE<�K�� ��&�sj	5Y��#3�'������dGk+���9�i�Vv���ˤu���!�I�N0B�$�:�3K�:g�tG�������#
@�_�����i6��ѹ�t]�����)���P���m^L��E}�rJrs��r�і�c����Ph�T�4���BRu�|������t��Gs��Mo��Cڻ&.�]�Z������ ����4���������0ݑ����*?T&K$��A��	���hF���S����:�	sR�)n��0����Nz�[t���B���V]��e�bt��X�냢�:5�q��G��a#��BB ��͈ZYG�?[m?��"�����AWDnn�^:$�c�Q��
E���6w%����	ۮ�Y�8�Hza1R�۰h����,����qU��>a����qA���R��������wjN��wpzH��aU3g����H�3ޞX�x������吻�4U������