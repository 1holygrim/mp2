XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����xi�Ő�Up2\9c)=ka�W�1^����,g-HCO}e��GA3�9~t�|4}P�%8�ʟ'����7��&�hc�Y�ΤSQ�/��zxm��	��((MqUϓu>�0��-�D�R�۾�,�x
��s�ٷ`�����ͪW��\��c'�%�c�m��i��8�m�P)����Zg�t1mz��M'O�li/�j�&�����[��l6��i�V��P�ejdui�*U��$�bZ��)����� &%X�(�`[]H� ��z��LTq'�.�/)ޯYpm�c�T7V͙T��c\��l[�����i��~�|�Z�a*�?�$_>AB��}l���A�p��i	
dTT���g#t�9'�:�g��N�;��G�_�2��@��d'�_����o���&�?�����hgnE�ę���g�eq�,|�̀���������t�{���`G��C1�KPGK9�	|K[8^�������&�J\�6�ֺ��Ob�F�Fܻ,E<9X)Lv��V�J�Wf��ik��M�v�$�Y�H��	��H&e�
'�
��)�$)����/��e���4�$�S�"Td�qʘ��FI��4�dh����eR}n�JW~?���}"_��:�.wp�:��,��̳X�4��6,�X�~���
�+_2zx�D��j%�)�6�N�,���~��҄:x�<���,q������u:�q�EEs����Y+j��EN(��q��.�kP��!�k��Y������X�Z�\�sP�އ�$XlxVHYEB    7ddb    1a30J�<�7U�b����B����<j2�q'�b�A��!U{_�;�d��J��9�
f-Խ<6>��ʺ����^�B�ѻ н�~�2x�ď�����>*����rg��"}2|�O�K���S^�7���o��0����M�6�5V��X�|Q������Ņ� 	\��$&�|P�cà�B���tZ���;=M�R? �Ɂ.Q=���<��۸9�S�������g��Oձ����F�:Ymۡ泿Z�1}�w����ұ�6���F�(����C�Ux�w�A��g	J��=�\D��7[���3XY�o����t��n[r��7�A���SН������,���ST�I��� ��٫��&r��1HM��fWu\�z�I��x�Qh�_8h���e�N�ʓ\��d�9�]�	��\�$57� ���5Qm"%���Ԗ[�3�ܥ�2�a��B�uSݹ>�}k�����tX:���9lcH@�����
L*�Z��m4�0�
*�-B��l9;�<l�;7$Fl�,,> ��0�;���Tgϓ��z^$+3��퀺Љ�yA�N��E�A�^�Y%�!-X^���s�!6L(������1��O$!�M�5���Ä�-[��D�T�J��d[�"#L֌��O���	K
]������?gK���ʏ��Xu���Ʈ�:��H���  �-��bAm�⛉�<9F��L�}=�f-u6E�ƏC(J����C���O���F,���t�w�_�k��"8�hɸM��[���x9֊A��j)��A]���[�"��ڸ5t_���
�ҢZ���=��)]Y�;|�z9�m�y:~"˥��v����������Lw�����ӯ�(a˕H/5G/I&xI8B��A���L#,iuv��,0�U�'L��y��"�Xk�Cu�B���Ť׀-�"�B� �z��A�����U�2���B��p�p�K/�קDqRn �`�4[�8!y .��8��O�B�#�3��6��CЙ�igh8Ш̞�q��U�zIp!��6�9��	�꿉|�=��c"H={e���q�?�`��L�w�@���@�(#��E�� ����<q����1o,>G��?�
 �ȍ�FMb��_$ߥ��4>ߎ����5�P�X���T��k��ab)�D �{-�[ �T�,����K6G���#�[`��������ӴBE���l�(&�R�_���[<2��,���jEh����<�Ǭ�pq�9D[�4�QҝƂb+2O���'��NCy;	O�w< 1T�/�l�f�3*YE�1�J�6���.x�@����+�`�#e'�o1���4a�|�����_m9�Y^B ��@��2�Kx�p�p&p}б��rQ+}ڸ��#_�bw3�x�	�'���D�v@���ϗ�`�s#tUn���LY�d�
�R��#�9�3vtTԫ;;�B�����cA�W��Ƕ�}�/yM�Gy]i5���� &�ۤ��Y�RP\rc쟽�����T����d�!"�^�3n:�e�8�����B�U~���ª�����sE+�DHΒZf%ٺ"'�����u�7����_'N��X�p����3T*�UElk�����d�R�E�w�\é�b�qE�׶���I9OKl��+(Ixv@�ך��.�(��W�J����v��U�*Iw��ˏ�S�ǳ��X�dȋ<�i����Չ�9Ŏ_"���#��7�W.���iB��QdSaB=7���k�Z'~�ǡ���u����j�W0XUʊ���	�48N��������j��Vn;�=0�s.��B	��-�<w�_��<��~z)�l��&Y�����J�r�&՟|������[�����]S�&���J���n"�
���$���)�C��ţu@UF��!�x$�k�c"�0L�-s�!{���]��XLmmZ\���Ԣ������ET�]� J��0`���Ws�;��`j�u�0
v��ok��S���Z_t�$�Tqz V�	�E"X����풀����VU!�Z��[�2d|OM��8�!��0=���Ճ�p��0�%t�g���!�e�q��F�f�� C�|#�r�ͬ"N+�or82�a��񖞫�Z�fGʇt��W��������7��������i@I[�m�y��0N_��w/�y����iX��Ȑ2͇��� �|�G�购�YT �"���=R����Bg.�<��KCP��g$�VW7�tÕ36��M�2S>��W���.*ր�T&���=��Y'.u8�\cβ��u�_�X���f_�������{����|q���Ʒ�`�0>�.���� O�i��E���|;���vt��W��8A��IA�)�ʿ�mZs9��Ŏm�RJ��?/��:������O���|����b߂��#H um��/d�d!����1� 2a<�\<�
s���ml����e멺��i��.�ē�9
W$�*��v5}��N�(�-[��IO@3G���@���2��`Z�˪�<�Z��TY�,-��fE�风���'<`�Ztk6�s�aR����<�^uo �{\0] p�S��&C8�<m(]-@6��z�,��P;=r�mW�4���.;i��h�I!t��uI RDDݵIC��^��L��;�o}"�	�S�w�����d�pP>�X��]��^TDL�I��{�y��80InMm='�|N�&��K��a������o ���#]�)L�������L��pó��" �s$'Lh��/K��l��"xi�{EO6�I.���/?����iZ�u9!�&Vd@��I����S)قh�)�_?��
�V#b�x¡����=Q�_�nvx�t�����0��?��$�&�˱}�Q^�U�����V�V)ɣQ�h�i�রu������)��U�"��AR˓�^�y���k�a�Cy��括l�)�%�HHt��. �*��w0
�ʃNZ�u��jiK<5��qAp�����z�������_�WT%�Z#��bh=�~��I���毩�%O(�e"\�>9�~���"ǀ��/�j�~���qڧ��/uSB��4X�O�y�A��x)Y�ɪ��|4�K�	�ߑ�NRI�I�h�*in��ǒ�Ta�%�V�idi	π��ϮZ���n �Ak�-?�ڏ�
�qܝ���iƝ�R��nXeQ�$Ν�?�~�r��m���u`h
	^ґ�J��:�~�"�B`F�J#/�-�qH��������g�,����]������FB�=l�ô�s�6XE��N�6��E
����7 Ѱ$,��� Vo�.����؍��W�<j�"Ju��-���O<����w�0&���١�㫎�tg�<��	�2�F���=zi �;WG�qp���~�\P_5WiZ�*}@8�4�0��|8βPO�kq��4���?u�}�o��'��qd����z<�{�F�4BW�M��Ǿn&�텢������ɗn�~U��N�Tb= �&���D�j�[�o��޳�F�i���ʖT_o�B[�Qg7�؏�����y��A\�~-!jvKUO,�q'���ؿ����X�b;�(�X('��c����anU�Adn
���q�3�����Vf�����(Z��=�Ѩ���sM��<2�^�xyQ䅢F�N1e��3�����t)�a�j�����|�w_�)���N� i�"aa|4ud9������D�D��x9�����o�B8�%��UkA�5�.�v���6�
Iu��0}�evw8vnܱPײfb��CR^h����P@\0.)�b��6BN�#�l�d��(#+���풬99v�K+-.`r%����YG���<.��dģ �Qv6X��,S��r徘p�L]k^$�y�@:sI(>;#E�ŀC�t>P�Χ�e��+m��?�W���P(�S֔�L��F�
.�t�����҃�엸Ȍ7�7��<QrF�V�;x�a�t��>Xw,9&\�)7͐U��$�胵	�Tl�uH~��:���Ӯ9gbr�pf
���Aeg����a�V��D���;-;xr /�~ܔi��6������ Z��ȇݮ�:����i���tm�n��Jd�	��HEOZ��g16e��H�\og���A�E��8��������Y �l�����Ȑ�X7� �����/���×!�/O��1O�tNP	J�ύ��eK�\�������<��:rQ��Q$p�!�Y�9��s!F7XƼ��>��S3���0FС<�O�H���l>-�c�fTk��|Y�L�A��Iؘl4���ԡ�GBu��T��Ӂ��k�ZYj��2t��}�7����Eh"\�MW�T� ��Ϸ��;�aB�Hc���`S\��ff}�%T��~�G[>���9�w�_�J�UR���rfi%�)׌8I�O?��� � �F���\ѕ�]��:����*���|BX����*��2���:�0D�6����'�˪G�Z_�E�b^(��/���/t2��v��P
�{rPdX�b$P�Ղ��b�3����26��f*��Kh8a2�7�+-�)��Z���S�.yَr��|VĢf%�Gc�Y���/��ݦ���D-�ʝ�O�s��[.�J���F��N�(pɝ���8�����������n�83Y��%��I�e�`ڤ˕-��q���0qxȩ^m�g����9�ˢ��$0��LH�}CSQM���3�����Ry�Kz]j�@�Z�b�3s�rg�y��I��EH�w�c��0�L"�ߍ++�xo���������2V&����+����>a��!�0Xy��ݾ�)d?A�;�˧��^��f<~!IT�v]ED黎���e��h'Z��^��&g�7-(�Dz*F���{�Y��o��U�>�a�,nv�xCǓQ���Q��&�!˕=���X�]�«64C��zNX�B4Ţg� �x�|B���$؁F��j�=Ω�*�`�P��U$�_	��j�@d�AmV�TuXʆ�8�e�*�Yv��)'����\��um��>ag�rr�����l��Fw*�����a(`�����K����`Þ��ߎ���L�l��	�,�D<�����#ߡ#���f7&��
�ˢѮd3ς_	Z��\�7���߶�BlD�*0�SV��u�`�#� ���O�������s�ޝ�/Re|�\l��u�*��)8�N��2�[gB.
�aj�·"4�pL�X�5)�U�17d�lz ��]�,���16m ؝�?���x��WF}	����#�À���bY�l��T+_}]��\2���)���a�6�6!k~Gꥴ3�=��EF��w�*�*Y��҃*����?|��_P:P)�R��+��Ĵ����������t���6�D>�\ �Һkj�j���zl	��1��m�d��G�����{>�g���9�b]~L9�S|��5�"(|k�4��rγG$e�-}��Z:�F��K��7%��fV �ϴ�D:�Y�+T&�=��YI,��*(>���Y�$�� U2x�s��!fo@8K�iiY�Zܮ[�UC�=b�'��j�د��g��
�	'��c�8�hj��V�o�;O�4ʻ�q���^�p	'�b����ǻ.�D�/�w��s���iͬ����x[of1B��Ђ��(S>�{șc���wT����,_�}�AT�u<����acK
 \nww"7$�n/�S�oX��B��w�T��*�Ҁ��ؘ��G��������]�0#��)���g��\2s����t�����u�ї��?NH�;���S�e������D��_kC	&Ī��(艟�Ҳ��p�*d�������������n]/�ջ.�s$-��A*�G˰lB{��~#?�H�p�<t��7�-�=��$b��>/�wT�W^AH&�ޮ��ļ��~TwφFE�GF��&X3��0P���&B�AgpG�~����iR����䮇[A��+�]���T!+��W���L�3�J�"�� �g��?{-o[A�ogr���@wN=5�p�LE|�{ęj��}[B��y�+@O��3�#ۍE�� �C���]���e�����)�[D��ȕN�v���1MB����5[r��(z��\��w�G*�<[q"u(|�i�Q�dC5i0�2�AzW�=�$���E�d܎gݑ��GBr�������T3�h�,t--�|F��RWe1�0k!��]���?�-Y�I�ߩ��#ؗ�w���
�F�˫�2���(KK���v�Q�`�E}L;FH._5%��I��xùE�b����	�q����J[�q�����r+�q��q�zY��6�k.�ˡX-="���	�~� 8�n{���앐D�X�[0{kvL�˟&�N �:_�"��v��:[�$��7�����g��^N���	x[�����b��@Q�YD���(]P����a���+�4=5��0&hJ7�7乊7,"#�-j�Rw�c�%B��E�M��,��yi��\\����P��ǌ˹#�k���/��S��b��/.z��hʗ^�Vw�fk ��M�rfX�o	c	f_ (7P1�'0ؐ.�ɠm1� � �Pg�
���ҳڰ��q�!S�H ����|