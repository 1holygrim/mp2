XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��'E_|���U'�hy������9�H�+A��Dc�2�P�A��G���k@�`Ճ�i��'n�g�B�}��W�9-���-$�K�*s~��2se@68����]��Y��+��Y��]�o�(���-"rr���Ҡ�uş�P��|��e�����p�q��KS�������o��X1��,x$���r��4q���`�J!RaP\(۫�|o5�3�ͽyJ�p>]�a#���4�y�CrbbW�3�q^�Z��<>��r�ڃ���s�2��\������})(b )�O˅���0����}�&:�ry�'�C:[P,�o7�,�\e��̼/�|]#<�v�b�����A�q}w�m���Az)���1�RS\rX57B��d��������).S��8��@�;T½s8^Ǧ��GU�=N#/��L�Q���}�@��J�9g�y���/IW��q�^N����+��'$:���^B�ի��R�[j�N^ـ�� i�H%��c@�� ��M@�:ȋ�"��wD���1�gdg",�b{�[�p�e�ƣ��쪛y�:e6�x�����T�&�?%���:�}���P�NPFp'�Kq�iv�5�����{	,��7��Z�:(�
���u���ᔢ�n��&X�S��հ�Z����4���P�/9a��1�Mbn�j	4��u�9��Z�g�H��BF2�ħ�ڼD�����o�қ�,+t�/���Ĳ���:O�#W:	�2���DMf�a�����d��XlxVHYEB    6653    10c0����J<F�v�Sb2��
��Z��Ar����o݉��Bv��L����:�K
�`�"�,
s����������P�=�`��~<���0� 7[#�W%�2M��&���k��N7�T<�����B@JD4s	�s>R�k���[s���A�D@��S�=�G�L�[����ݧ}�T*G���D���}�Ho���| Z���UՈ!�AVv��p]��8f�o���Mlu���u!:]ڻ�@zE�AI�*Z7`��#�G!z�����bb�D�,�]0��&��\�׀�����gI����22�/�G[�@���`]�BTTB�w�g|�ٺ���?�Q�K�߹��W<�����#�D�.�D���-�F�<���T���w%���ʮ��XoL����)�� ���ĳ��Јǻ]�'�H�FY��ӘV�HI�����@����ש�-�fr=��.�m�S�yvuBR�2e^�puM\(�V�x?��l�g�k��0�l{��\恈� �g���s�7_G�`M$h�����Ȟ��K�A5�[rޖ�f4K����1r��[�NM<�\։W%`:Ѐ1>J̯�����=�AHGQkԘ�eo�����/�a]��3c�	R��8c��7��_&���_M�<��ồ�W��S�&��!J�}Vٱ�lG�7�(S�Q�'̙5� �U�vP��b�CSط��ZNPf��[|�+�ӌ�������LU�@�7ť��Ŏ�c.�e��e�^$la��m�vg9MB7[��������Y=��!�e�*Bڑ	y �c��qL�v��9r�V��>sW�F���z[����\?�\q��;��<��o���Z��u+}�@3C�H����w\OK����,ҸyP�!��>Q]�[�1��!,D�HO��W�G��N �lp�4|�pޞ�J�zDN���'�����u��Y>SG*!�u��r7�󰭑A9VH�'���`r ���X_J�4?��f�4�4��<b�O��r�?�M:�JRf@*�ຂ�k������I�],H��ʙ/�x߿�l��p'>nW6;a��F�+O��u�9,�=��~�C���7
8�P�z0��h:0}�t 3>�?#�	��A,�9���{�߫�!r��x�=:qE�׏�a��U19i[خ��ψ� ܽ��݆��������N��5f��Q�G�ªÝ��@��'D�4ն�포����"�(E���u����j�s�B7�����l�K3�s�_�xh��"�0!r��`T{7�e��k(�ɅQD��rH���53�>Y �A�ި��+G�~'�YvAK1~"�d#露d2��t+���,m���M�s�~M�M̵��F ���r����n.���nV�ru�Vm��GG���������}�l�����v�G��np's�}�������!�a��s�Vf*�
�_Y͂*���v3*����LHx�D��Rt��L(��L�����k]��H�Vl>���k`Ը�T����|p)OѿGpD�)���.�[���|D���[�p,���6�|�jקїI{���D=�\���%�*Y���� ��!%(�J�X<%�b:!׿֤���.���7mq'ƶ�Kw�}����m�� SF
�9&P6� �?�hFv�p���н�����T�
��Vr6R�Żƃ�@:�h�(�Q@��U8k1�S&��a 'n~\��8ӈ>"�(1��,=��̆z�W�J׍
_�c���[5�l ���Pt ��grq��@�쌑n2>��t�b�%��-}�!��,�T���3.�ᡤgǻ�����W���F��u�0�����K��'_#M���T-�r��#��G�X0�ոy��j�)e�[m�4dq�	Y�է���{��s��({����5̆e>'�v��u#������"?[	�[�9�*]t ���Z�p�n��ׁs[u�xJF�.��X}r)G1$x�Zh��c���FIrW��zV�3d�ӊs�oE�U�9N��P�)�������Y�P�0�������!83����Y;��Y�t�iyI�_;s�`��܃v��Q���9�O	53<K#Hy�d]��ad��w)A���;�D,��*�3�7�Yo4�+�n5?�����ྮt,V���PK�~��5c����{E#��.��E5�&QN{!.yTA/.֯�����m�|}��{ꋞ��d�]HZ�lT�up�V
�l��֭�6aՠ^��Y�å-���+���s>�+ʆ�2�O�Q�T��rШ�:0�$�!,�0?��0��t:$��y�ZN�.Ԭ2hP��%Tm�i�w/��E%��(L�P	:��_ډ�ʉ������P��B�]B.�I@�Y8��)�X`�$��G��=ժ�����x�U���5뮩���Z݌���m#�,��O�� ����Fas�+�a�N!$�@���3�?ZCb����3ꐹ���0:��Sr<�!׌M��P=�1��B�%w4&�C)��]�)Z	I�
�8���¥�t����J� ��J� s�xK=����<����=���_]�!�>U���'zH�4nl��{RӍ(���Cv���>=��R8��(��'z^6������<�5OTYE�h�4s>�B���j�s�ЁN�u�JQ^hR�Գ�T��I�-�K�D*���Y�F씠r{64.����@p��V��$��Yq�ƚ���
J~��xy���Ժ�W�V���wKeP;�Ҥv^_�� ���Xt��r�YzC�<S���{j;��$���0^hNHɊ���K�1��=Q�9�|;��R�P:o���=��)`k����9@�EE;K;��J�g���id'1�j���Y��Yq����|U���`v|Mx��A,ݯy\(D_��E��qSb�~#�a�b�ْ�ӌx�:i �2��e��|�ڣHY����ۺO��W��uLp�C��v��.�Y�Ǧn�ѥ���Iw�f�,,�V�?T`Պ]�əBGi�ն8U�]�z�c7G��~��UEL��O�?��Au��>I(ҁ�r���N�%�g$�M�a��]<1lz�W���	kXf��.�V��_��49���p'4���P�%#4��]imʗ�s��h�j��8����G�@�p�>}�D崉/�J
�g�NU9C<c�����]Y�3/������(���-`��Fù��N��U�~k�lr5���4;�T���\\���� ���Ns&b�z�h��r�C1�3��3PmЂ\�S)n+����0c)��i��$�Sܔ�ِ���0��'ޱ��Kº��`��d ĩs���=(=P4��(��RS���E�M��jaZ��ƃ/������� ��|K,��������9���N�麗ê����4Sn��M��yJn\�s��6U�(�����.�
>��Ln����)�YYc���3j[[��������ֻ�^B���=���B�\؋��h�Z�:�j��}�~�i�d���T�������k�~�����x�ܞ�sN+>GF�:���o������GPa8"��jIċS|/�E��9Z����+x�%�@\�}%���k7�w\v��0/S�
&�NQr.ΔS���]w};oZ�W�Q�����~�	�JoZ��Jf��~���p���������2�챋����9�Cʻ�J��~�  )��z��&�*g]��_��.�S�.Ū�����.�iW�_�����pR���:�X>e��3����/��p��TV��PVݳb�FV�aR&|��|OD��ŷ�ك�a!�jj��s�س�6�́�6,��t"Ok9��V�@-��\�\((Xo������%�#���\L�۩�ZL�@L ��pu�)���-��|�)X��J��a��h��(�ըb�O��d����u�����;۴�]c� ��)�� Y�_$1�"bQ�B�V�����;�R���t�IE�l)�}�2�>���WQ�UK��ͬZ�^x��lm���DJ4\朇1�~��� r��C�]�V-�T,�D8�,;��(�����@�_�a� �ڂ;w��L�Tg��_�[H�&^��"Խ��������u+Yu�Ea8��=wݑ�X��>T�+M�S����	d�����<V��~��dX=�A
�E�,��G��r�2���Z�M �C
�dU}�g}f��\����P����v��k%S����=o�G�M�