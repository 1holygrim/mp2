XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��o�|�P=��`�	�4\�@���yA{48]������b����|�5�(/g� c���=d���,��$�F�[(��J#�&Xw��G�Tt�JN6�m~����$a1��)KW��Nd�翍� �:G;�`�����V4@���N��=��>#��"�'�*c,h�67�`�;���g�XZ�ۦ��R�6N���`V&SV<����K�?��$5N��E�T�S����"��E1��Ϫ)|��H�\�Y��6ߊD?*)��n�W4�|@CDvb��sǻ�+o,G}�47e{���zM�R���a�l��A$�9�R��oG������\ ן�֢pU�|��r����z2o}u=�}AC�
dl�O���,��,�Nך���@y8���O��屫�`}�oa�Ƃ�g�&A�1�Er��N��E��`�q��}�~�e�$���=�rאe�(_�$�(�QJŎ����G)$���*�H�)�䱖��Jt�@��2�u�0���-Y�}�@�	�r#�i7�]T�m��b�@�q�%��U�=2�Ȭ�)����<ˮo�ӎݔeb2.��%Ы���S���^��"p��fw/S��ư�L�0f�<ihl�;]�¾c�~{9":m,�(��A��-���ظr朷G΀0<��d�'��3m��w& �M�A����8��0��Tmt� �+�e2�#撌��l�{iy�\�N�H���M+�E^�N���m8}j哈�W�H	�W�E):�D�c�o��Rx�ο���XlxVHYEB    a0ac    1e80A]�4kc%.�meӜG���$�;�)<���e,�DK��G
�)(�|�߷�E�6�0�C}�m���������#d���� �tD:Wp�8W��\}����d���l7�]�4ao������h�`	q��� 5%�y����fE�AR�Y�*Q����pP�3�N�s����p���̗<ʴ���f9��F�}:{����U�P��sseWۉ�v09�c�\��?��&��@��m6�¯��瞗���L;n�xb�k�䑢����U8���(��g�ͳkhگ�(	R��ڶ�ME񅶠����͚��GJ�}HlE��,�92�%�D�7L�(���4RXh��M��&�ey����XA4���FJi�'����I�Ӯhw?�b�~�8ږ�?8Pt*��p~U�r|���\��uw�{2���Ԗ�5
�Ga� ]V�������&w�Q��.L.��^�^����{�&I���YnYO��Qb'!_0��}�̛����|l�e��Pj��-��!�+��vf.V�ݶ|娷r���(R[ ��{�Z�_�r�+\� �!��˴:��c\��~�葌�t k�[V��ijD�F��>9��a|���/!�X��>�"����%��
�.mf�3`��R1$�cn�0�j��d_�x�dbM�G���!�	Y�ָOJ.\�Y�� ���Tؗ��;���Kd����ޑX꒷6�+�;���`6���������V��-��
m/���C�*�j-�Z�������������������Mw�{)x�
�~�e�c�́�m��C3s�uu��l�|��Y����Cυ͔]e -G��N��R�$s҂�X�g⚗�dR�@�Q�#�èw��S�#�.9�]�v	Q5A�j�]z�*�L����uzj��q�D�?'"a�V�5�nI�i�@W���?�uh�(��*�E`�k�/�V��|��H�|�6��p����D�c�{tU�%iҌ�i%��~$B
c�}�e�-��^9@4�����0[DC�)Xb\2V��M��T�F��T��^���H��q�~�(�q8gC��B_�	e<!�'�ʔ����b�ח?�����}T����;�Ga�"�p�B��_d?w)'�(�^`I�I�W\0�H��kb��WC���^a�`1u+Yr��$��Q�P9�Z|�H���Z_}�� �_�"������C�-C,ܝYo������w�i���*��-��sC�`���|	�M�����"Q�GMa�{���7���m|�n�0X�5�A��3��Bn�]{�L�!`ƌ���sJ��'�s���K�`}��g��2��(77U���d�%sN7�(:r�*��fn��>�����lD�4�8!���y��%E�X��9<�����lT�)�hp�8�q��>��'��'��!k ��&t��%�D�⥣�rV9�t�ߤ�vr��-uBI|�v�!��+ZS��+�28�K�y�Ĝ�X|,�����W�ܝ"�:*o�ko"�_�v;�ԳX���H�Sb\`��T!V�\a�0��"�X0��n�u�Ȩ,���\�Gn��cs)e�Iv]��0�7���G���j64��-[�Yq�ǶPׅ�|��)�K�U���ͭ�邳�AD�#�b:3Nb�{(Z�J�t�!!������w]h��a�}�/�^9�����w ��P�䴳�e~[�����y
_�3A]Q*� r���_��~��0����sye癪gp����]��S���X�M6��U	��"�Q]?)z��2�ʋ�vZ7��-!W�ڬI����r����$_roxo��&�l#������	�^�<?jTe�Ζ��?6uC�d��� Sc� ��9ꔙ�ݪ�
��[�d�}X����N��_��qy�YcЭ<(�c������kL��HXc�QT*I;�H��Das�5����7�鹿<]��A�vp $�/Ţ�����	`�2�g�{��R����hOP��������y�����N��v��2�Lg����x��v�L�q��Mгn�d=�����?�iJ�e �[Ͱ[�!�\ͯ����S��E�4nVM
�A�%�~"���� '�C���m�E�b���8z��/������re���-�F�VS9	�
Y8���5���^j� ��v
Y����g^�;��E^c���M𾮡���K��õb焸Gfv��x��������&���v�����w�jQj/֭���֯\�
"��6���2z �.��aա��I��6��U>F?`�w�l�����aj�L,ssu��>�p �� ��/��*��UW��27h����S���|(?�����xe��Ig�6!X����~hGh���Q�-��K��,��oL
qd�j8Xu%~e��s�/�t)?���YoN<��D��Q�`r����VB�Z�aF��I夓�Z����b�Q����!��VZ�h!����0Z�,��ːL4ly;�"u[~��~U��v�|f��ua�'�}����L��w����B���压��Q(�(��B���'����I?,I���3�-DU0W�M�h�r�{�x����fXn<�H5���u�<EK��`�ȧ�3�l�H$�2$6,*ߩ��J���8p4�4s���i�S�a�� ��{{m�����(�V���7��i��5*�7�4�%�O32�G˵&�rS�F&kSW�����M��3F��X.:�X�cI h���/�>1�ɉ��z�H:s��Y.@�9����?h�C�3!~V\v��Jz���_=E��]�$u�6�CL'<����Z#={ >]z!3B�
"J�+H��L��w�Py3���C��$��O�l�^�'wۧ�-� P$��3چ���/�TS�����X�C�W6���n�\IR� �G����I��游��㣗 Hfu0N�vl��Sm�`D�M����ۃ��)�
2�L 6g���R���a֔^nXjL��h@�bc��x��|�pt��Zbk
���)>2�Oz���=$5z��!��a�ND=T"���u�z�;�B>yW�;���{ֈ',�xX�9/�r�h�:C֐�^��4tϊ{�'&��\�n�]���.тv�:GM *e���hi����ͼϹ�Sĩ���v�8e�	c�xu5])�
�𗛷�c������z�&I�pW��S?7���vq�\̽ku����>G�E� �m�yf�U���l�����ͱ3f����+��(8?�s�_kvBa���)ʿ�ch<�Z��[Պ-���-��J%Ij�Z_6{M��<.g���ة[�Mo����V�!���%Ma3�8����'����U������X	�5�j� ��v��X��q�}�s^�#`�s_`~,��裸?E+qR߂��a2nfâңM���c�����fb�jv�w�E�2up���ϸ���*�\��hVY�.*KxlQǫ#0Wm�t��PoW��y|��B��[��ُNM:�+t�G�gG�-f��0/��ҋm`�"��"ӌ�7�r��:d  ����j�l�Zf?Q�:�T�y�b=UȜ~\-�$�����ɲ�6Y��f��+��fhgJ[������Üy���ĩ��]�vw5,��|����+��)�?(21��co�
Na�1~������l�w�˜M#|�
z0W^I\m��|7�ܶy�A����P������g9��l]��!��C�-�C�+2{-�t7�I�#�Nm�}Mɼ��9C�ȿC#f�U6��������n۵�?�1� y���kV �HNH]	 ��J�^E]]�E���![iz�޷�����b����߃D��BR�!�G�3�r.a̙�v��%n��a&�=
!�J�ʀ�d�_?���O�B,��׽�.Qk����YT-�w�c|
�U�R�S�)rC3;��;�+f�����o��'	��$6Y ���Ԩ�u�քW�He�S���f�L(�l{�Y�]�f�C��5�<=V*��t~5F&�Aq���38H��>q�dN),m����>d�=9n��J�{����HN��_90�㐮z����p�W+\c�o�J��*����C+Fe����=����&.Q�ۊ9����aq�| �2��?��Fƕ�Ƀ��q*U$#"O�	q-r0$��8C�\cz�:�*�Io��%�F� �R^خ��ZtXS�-��f�� -xt:���z�ꝡ�V��Y®�w��OX��׏3��+>��v��M�,/(b��(�Tw7tT;�O�����ȥ�Bj����KR�k@����������]��~R��K��n���8DS�U�Ug,����mo�͗��o�f�:�$��	�*�ȴ������+�3;��}mǢ|���S��!pl�3����|�x>���²�6�tBSn�[j]�)e����1���|�vJ��$� ��ԗǇ����8��zӄ��I�;Q�@���f0a""�MBAͻ�w~�U�/�`�iqmBv�SJ5�#�Ŷ�	m��u�+�����Vw�NYӔ��f[U㔐-S8Br�&�)�w�)��@��q�px|߯߃���"�:)�����������E�t�UY�L����=ֺNbZ�8�-?L���'>Lm
�����i��\h����6�L,����8���uZ�QZW����Ygtƨi�8:8�Mc������n��=z�)������H���i�	��T� �:�����:T��p5��R���R�/3m��l�X������hou����/$�׎�4��n�4䛵�eO���*�a}E���@�2C~��G�?D\��2*Qf
���~D�KC� &>I��h����Yz�!L�Kն��Xe'�&C��k��h�=v2��
n�f�Q�o@�����a���N N%��!������^�٤pHik�ؘ:���i�^���o��pɸl���aߠ̭z:�R�yqo��"��	��D6N�I��
�*%�u��dd[�hG�.~`bl�NT��k����7|�Q���<f^V%V����$*���>�'�p`�!l�d�:ҖWGanoヮ���'��TUx@( �_����(Z��xE�K��k�tais����P�Z��&_�ic�7e/��� ��ƴBgqQ�u�>���![����[&B4��MV�����?����<�[�![�>���+��S3.%�n������@RUX|��z�q%e��%�Un�����:��X}��[���ky�`�g6�������j�<�����Ώ�]5��JLg}T���ߡ�Ȩ(:@����p"OP���?����e���P�hF���#��� ��N�E�g�9�����K~D���7nz�F4W�޲z����Nw�}zF������SEf�����_v�������hul/����7D��sH��Q�̴{�v�V�5&��T��֍�?A�ξ��X�Ļ?ͮ�K�ˣe��	X�Ew/����s�Z/[v�b���<�"=6�۔� �O����"v7��+�럘�����/�<��ef�-'���ˏH�~���CǢ�J�|����5��%��~�B$8W��.��J����M��5� SY]�õ[s�L
�/�Ң�;�l�Ir	��{�Z��,���͹wdz��zLOĉQl���bDQ"ʾ��q���s�S��ٶI��m
����m� �@�y	;��'�]�4{[,�Vk��7Z<4��p���9�������a�Z��炱Xz D��ut��ȕ��'������s��N��_]]����͋7�0��H�E�.����E9(���3e۶�����E	F�S�Ö.A���3���X"uD�O�j�?�[pU����'|�М�=s�ؐ�ɉ��KUd ��)�����_��K��H�0�I���tQ{w�/�̊���z��f�n�?
,��JO4�\���Jڎ�O�����L�~�m��<��{n���V�`r���������Δ�4��E�i�P�88t��DuB��jHW��&!�h���~�suWl�OgNOo�v��s����0���9��0 �e�E!<�(�$>���\�w�,��9lU�;��<k�b°�Y�5eչ�0p�
���ۢO�N�v���Zp\-��.V�Kט�׍w�ojY��~�	Ȣ0���R�������x�@X�ey��ty�|��3< 9M˽��Q��{�����}±a6����ڮ��0 �(�oJt@ 4Ù�J�����q���]VE� g$J�s��	�\���GS�G�.��n!ՃV� (}H�N},��G�ȕ�a4�QP&W�7>��AN~s���ؿi`���	�i{����Z�n���C7��_���nid~�@=��q8-EFm�0	ʡf��Ń�)U�ɑH��Ŏ'd�T�6S௃���t����X|�6(�`�}��}@Ƣ����Ѩ�8������쪂Q8���9t��ֈA�hQٓ���=�'A��:�*X?gրZ�_P;Zd4I��bY����G�O1�����x	��B+�WaÂDu.B��_Egi���.� qKw@�}p[>[��<PM�������A��mq�F�7����ч$*���i�sb�mopa���h�Q����4>7�U?�Mn� a�*{΃!D�0a`p{�������͕��]ě;�9�㚬JH���Zr�7Υi�`�,�D[�p\?�L��mI�����t�U�NH���	=�n6�) Ȏx�+,5�3)"Q��EC�r;s4Iǥ6C���T��_bS7%/��72�Μ���{ƚx)`��e@E9����<��S��C�y�(�^]��nTA*:b\�=���	`ە,)�@Lܕ�JW���!H�Ie�*M���ܷͬkr���U�� ��b�	�5�P���@�Yއ;\��a7/T�3L���(�js������K���L�v��J��� sh�JM�uZ��f���N�M�@�"�����7J�k���\`�75��j�}}]��B愈<1�73V�BY���ԟ�/Ď�����,	��6�X<F�F�3���}�Y��2|%�:j;R[�D�:�9��*e3\�G.�昿���� :T	Q9�O�y��J�N}���vrEַ�s|oy�_x��R��B�1<>�
�G��m���mNh�9�.�N��E���F�{�$P�@�t��*1ϩ$ɽ�R'��Y�UW��b����J���<r2��j^�(�6��JG<u�"x�_6!H��\y�i��u&���gB����S�x�Y��C�c`�V��\u�ʽ��;Y:uS�=�`Ŋ���B��.�֍�&eD/}���Q&P����ќ�?uȨ�$Ww�Ҕ����@��_au<+Dj����UT�}A%`��S_M�h0*���Q}�����&u�X϶��3g�)�*W0�Wx�+�}�G�ȩ讐z�m������_������f�%�e��G�����W8���)q@�U���Tx0��z}D�	 �0F/�&�:H;�����m0TXp�"֠h����wW����e�Å��$0n�|I�M���T镴Q1�v]m����fyN��A�����7�H�o�:G�l�ы���A�������7�C7(�˺s<�����\�\v4�P���#�|ih)�g�d{�鱗�JW��d౺\�qp^���'�xs��/�T���63�2�y&t����z�e�(P����}8��b�}dvO����i!P7}]ӕ��q-V����*��m@k�(