XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����lMr��'y,k�t��z\`���f�>�3��V}���j���7#D�͂��s'�TB(5��\`�"��vc��_�l͏�*��ޅFJ?9��mWdz�h�qt��m:���s�$���q�ЈDa���~�N��-��S�)5�qW.�q8����9L��J�r�q/C�d�����-�x��;8R����\L$��)�酩�!x�}x�t���p>)�����(sXj?�̐.d�����\����#���׵8x�Ȟ���n���֝��M�q���Jr���}Bȶ�ad}`zp?���a��
�Ƣh�,��
2x0r�g�\�=S����%l���pwݘw�P�.�ďg��g?��SW+��Uhր��.J<�k�#X�q�����#��}��SZv0u����;���&6�K�'C��AqZR�W@k���T�L��i�%�^`,&��	R�`?\,��y��Ѡc��B��(7�'��he���1ۻ3� م w���C��.<��eۖ���ͮ\'�.��>�7�+�=Z5��>���=�Cr�7Kީ�� -��l �u�e�l�T��3g�'�����uy��HMd~��|�����v�:l,�厽�Rty����_I*�e�B��1���T�	t�n�V��YG(�0'�Wqr�VI��>s�*��A�>�W�ˊ�
"s��_�ggً���ʃ�����\b�����]�d	�t���������~K��g:'�����`��hj�p� ���Ɓ5NXlxVHYEB    fa00    23d0��8oY���`�.��%��Q4Ls�N��Z�D!Е?m-}���	1�ۄc��8&������g]%�E���au�<���ޏ��;�m.�e��\Z�@�S��a����~9�4�^txp�q�����:���?Y�9����,P~��$�������*'��_ViH}�3��y#y��>��K�_�-k��AvޚO�RO��P��Ҕ\�����\͝~e�x/����c?:��x�\O w*d��]K@m��Rrq����ftg�.��,T˹���D��.9��%�".�Q��
`l6D��>�ÔaM�z��������]�uR/���@�I�R��r��a�,M�D��M�G}��2,��ٿ2�{Hy�dp]�U�(�C�Ռ��AU�t����N߫�墢m�d,-���)�0��C����t,Ü�y�L,y,*|	BE�Up%�}�Ӿi�����p�|�OqG��/s�ՙ�`�
�e�Ó�~��vrL���8v��y����[AٔϠ�Bt����㋦��A��DP���9�H�8u�w.�AM�p_b1��I"��4g����:1\�!d0���0&
�7Sg�ǗwU�]��bb�m�e&b�Ş؛IO���T�xCL>^���1p�.▖~k��M��h?�@#T��:W�e� }�´-@����\�^��L�̹�p�<�ݙ�ہ��~.|���8%�C���S����\Y��I)Y��I8�҂.��#�0p�Y�w�(lm\��F�7R
����8�y>n�>�]���H�A%�e�������{67[�
򻃢��X��)�����ؚ������R�*@E�dn��7?s�,Κ��r�1t�ğ��~���6��q=5��C%ߩ[
��#��mT��Ȉ�G���fQ������f'��D_58MV�����/�-����w���ǣ�;�o`� /8C�а= � )`+�8\SCTp�\�Î��'����j�U�^°Y4��/��-�{��c�T�U�c���4l�Gt�k�
���LRjM8���<�AP[���=�F袤�w<͝6]QBhj�&���2�����0���ˠAXU�RW�� P�+�X1�X��7�MC�0���ň�U�_�ZO�5��&ԧ5����Sp���]���ԛ�?��,Fu�0���JB���u��l�3����仛K>n����o�.vl��DG�8g�6��D��͗���9�L��TW��f��#`%j��q}�'O��6��v�*�n�on<�C3�Ф�/��ՋN��e����D�{�=�IH29�Ko���\�y�Ue��g���2�.3�0A��q�o�aqğ�/���!Y�%��OH�o	��(�7���T�&���8y��f\�0p�g��_7�]]�t���CW�t�Wl*8(,�s�:������G�'}��c�`���4\=�S���NۼF���[LP�f���6|�%'VX��h�/�K�P|�N�����	�R�jv���ӴQ3J�ţ��orټ�`R�U��gt@d�T�-�Q�F�R�o��2�0WB���I]�rL�dic�m>Z����2ܧ�y����Kr!�A��q�6�M����㇡0���Q|�W@	ShB�O�?ώ���m�<-��}l��4Y]atA[-ka�|�?��b�*����Ⱥx�H�$��+��?	h��`�VQ���͎�?V��]�>���������X/�tb�;f~~�F����2��|Oe�w��%)��Ŝrm�$�1��-d���11�r0)�����o?U�F~rd�'P��I�B���l*#� �vnx�A�$X'�(���AF�ptu^є��Ml���>����N�-�d�������t�B� �7�$�n�,}�]o��,h2}죷���F��O^����D��:+�~>yr0ihL�����zN�������^'�'HQT:���
	P���#�聭M���`��҈�r��g�Z���<��#�Q�0A�'4���N���MdW%=l�,�rP��O椬e3#�$8TXr�$E��`㞄f�QF�{8<���?��a	��5�(e��x�.�E��o��q��2��Y���7X��fn�9��>-�����_���(uk��Ǻ5��T?&��:8ݯt��=8C�:S�@�(��[���&�5Ǟ��q�̡�CP2�O!/���b~����/ �m+��y��#[N�Uv�.�*���]��s���)|w��%��H<��dYb�0^����D��q?�� �W��Ep��1ɯ�{�b���/4j�6^��� �Q� {a���������h���3�� =��VMR�|�HJx���Φ�a��=M�)�,w���0����)�ڑ�W5�e�zu6����Zj/DP7���zN�0��7�E�*�wH�°6���wP��/fq���ݗ�_30X�#Z�=B����1�>ׄ2-[��*�	_��ީ�N�_[M��\���F���F�B���Uw4a��$��T�v5��j+�=���Ջ�w%��A�@��e�q���./1�-R���f���dÁI��o�YOo���ؘ�H���t�%*Qɽ����U"�-wL��Y_B[��F����F�~�(>����[5�Y��a�������M��P��C55 ��՛�f�0�y͒�@%�ԨL�s����)������ժ��~����N��L��yP�� ޜ���7�8����ʱ�Ԃ�?e�F��7���tZ2Y2�����io�A����Vo��d�γ��$X�|_	��B�왖{򜆫�_��WS�z��	��ˏ"�x��)�}�%.As#�-����"��'BiVYxg�y�Ϙ$��J �����{*N�|�vi���qeH����y��y�{�5G���LI� ��/��c>�=w���W#Z!QMগ/h�pn8�E�E�� (����;=�iF��B�J�c�υ�����b4~�EjPZ��h����(xg�V���p���q�od�����Q0�	�Ӡ?|ҳ^4��b9��X����4=�M��>�\��;\�B�8Wf`�'��yI�#���P��{d���$�pp�{�YK:���	&��D�R
e�ۭ2?���K}Qr��cr̰z�|"yE��'�����Hش*|Մ���쇼�(�|��op�&a��RD��%�l�vq<o�t*z�³�p܀yDVĹ�$}�^�,�7��v�T �f|�($8�p�$@��������o�Zf()�u���Sp���"CՐ,
ᑔ�B��Ie��<%>G�u)�rF�L�7���TҰ�^pD:�/��1�R`�_[�'�_�M�v>�&��9uw3��esF�N{�����ڛg,�;ݧO�7^�$D��$��������	�_��Or��e�T�&�s%Fŵs�k��P!�K/碦�����_��jD¤�7v�T�����iC/��`�l���dI��d�\�!��A��&�l�����,(u`�Q؍�"����:QuEG���r��������u�\�/~�_��g����R��~�Z��}D�i��G�MCݬ����\H��M�#�#W��׻Os#p��3��*���$������v�8�n�)��3D_��d��b�����4��ޫ-�c������G���Ȏ�R�ڣ(z#� o9�W��t?��Ր-D�ymbmT��7��l�#�
E!+=�H�}<��v�n�ԈS���I@ʟEIж��-� ���f���f����̧c�!����WJ� �����e8tE���Ʈ0}9H!2_�;���������'�Y����E/㘕�i�v�-*EnM���I�)�a�^;e��I��\��˵�]\�텱H�x;�X��U�W�7؇��i:���~��=$z�x�U;�J^�ƈf��C^	�v�5.u%��dt�2�H������)+7�u�b�����\�*��!%���&4������JNv���>��/�P%%�,i��A�sܫ\꤆���������})�9���='��ֽB=��.��1T����[��I*!s})���,v'C���[]
{�N�dg)u�s\��T�4!��>�T�{�G���zC����tj]N<�;��|Xz�Z]�{��|RL���b�J;����z{*��D�
�`�#��Gy}ïB��u1
�\&G&�pJ�(���"(��*�S*5YG�*h_����
w��(a������#���>Oi�Z눾#|��=s����'���St�b�A`	? �o�R�>�"q{@�-|��s4n����v5��asC�7P2�L��\��Si�k���Sh�����%�Z�[<���W5��������Ւ�� X��㫮L_�2oV���py�F�0�e?��`��^+��4Řૐ�2��ï_��|�y�B0�Thw�:� #c��)���I6�1twf�/�(|����@p� ���GIf!%��*�9��c遄���n�Y�~锢��-�2����_���a$6�d��nm=���/p/�t0'A�+�o�w:�6�Y)��S\���y�
�ba�,�Sq/��������38ɪk5a���bv?�aP�f��?�[��j�rI�Z��.�$���$/��d�^�7���
��V!�+���b<�JJ�hx2��D �:���R�!��T7�K�pCf�)��Y��+�Q�1ڱ�����v�6�,�dԣ�x������Z��m� E� �LG�#3����=�x��8^���1�E��vȴ���!�e�/d���׷6e(�̕)q-��
���{�j��]:�1��s��I�F:�Ev�}I�L9Bc-V��U&:�콻��s�9=��d���qʛP�������Xޗ�n@H���~-����E��|��R>Z%U�j�}�qO�����w,�yub��p���,�L]9~#�������+
�#�u]�"`B�ڂ:��E�r�������g�tYtU��.���w㮟�e�Jk��g��t�x���}"�죚�!Y��(�MuwA��ʐN���N�	�Ɛ̆���2:�5�9�($��&�)2� =M�=A�2S�-#GT���ǂ�Z��v���P���_`�^���˱���a��3k�η��@H;��͕�lrn ��T^�W(��*x�ݪS��ƻ$������I������)1�K���Y'<���v��5HV�slv	�(\jF��b���1h���h��=d΂�j���U?���L�Nۚy�̝���7o���U)l2 z�С�����}����O�����E?E)��yE����ʨ��2i@�L��������?6 0:e��\_�;�rz�Wq*�n�;���������݊��e%ʘ�1/{����P/d�d�S[�,���p3)�̫S��u��L����q�D�mnk�H!��iO�q �#耙+�)�)hq�`4��_����������/�kC�B[|�K��*��5� E�c����9�#�z�J�j0�J�A��E��u�?1[<6���(���!�#v������i�;�+ >j�舗O>1��0��5М���Wi���!����¬��E�e��$�A�z��Lir���,�� ����j�9����b�g:w8�����8(Ä*~8�r�	�z�mKG�tN[^�(�]��'�T�i%�4�_t*Ϝ!�d��7��؊�y >�Y���L�֥�Q�-;ove*�� ���9W,�h��Vg�����^4C��e5,�6�W��%B���������h*5V�d�l���h�sɒ�?�nyf���V��`i�Ag3?�Ϊ!�q���������q��;���"��{1gy�*�4:G�Y2���&a������m�=05�ϖ�{�(ct�-�?�
B}�	�[��>	��b�Pv+d����Oֿ�!#A��)�&����Ξ�����g!y�9F���nE߯0z��Y)�㳝#����L�JJP_��P�A	Z��<�+��^�eݵ�f��ɴ����oS*;<�;DN��H�A:�����3ru�O������,M�Ȍ�����f��*K�bX��"�������
4�Lŀ�wT0j�)N�.8��r�j�ؓs��[kU}��iڅ�����&�X]Zd%x=�VǠ%<�H�o�(L���i?�+��b�PH0,�*�9��Y�g�灡?�ty����}J�[K�*��$��e+U� 3;ꉆ�����Q���{_e,���R[��]��wυ=�δz w�2����#O�E�n�����T�<�J$�ȭ�Z�����2���Z���mNh�Ҍn30�d;n��#�'~�'(_��N�Բ��(�%8/'�7/��)4![�,�Mw���S;�D5��F��x
�.�@=jlv\|�������0���(T�Q]�X@@�y�o��R��{}Y�M�V �3VF��pd�Pf4�3�9��ʰV���&���Z��_�HA�W�=ձ��3���tP���u�l��ݯyf��{���#b7�����^:ɘ���+��m��7䌱}:V��yϣx������ՕN4Ge?�D�h�ȇU�H!�X�&�����{�Ob�p����MfB�|Ҵ��u�H˃���� l��+b=N�"�H �&���Y�y�<�ؽ-���X���m\X�+T��.)#��%�J������T�_�xx6��&���1����K��4�p��q��ι_G)�
9��{�xW���LB䗲i�;�Ѣ�"�|@tg_ᒇq-DY�.����S�V��t��~�nn�E�a$����`&����SF��j�o�.@������?+�[����R<*�l��2�q�b�~��jtqQ}}�zh���2�˒���#{��{�ۥ��([�։_�ķ�2;�j�d�Z�{�BC	v&�K`�!�����v�c��w��������ż��T�	f�m���i��}�vVC��@�� ]���4��|��=؃oE}	R��y��8��]���;�̅@�a�u{����˛���E�$�\?�T�ɽ\�4A��rs'�C���uo��7	��,�=*�o#w���ʁuW���&���IK���B��q�g̅�e���fSETu��¢�9���[�]НE���^��]��|��:��L�v6l���g�?4�� �u&���899pf���/�,^�K�S�C��@����kLoI` s`8�@�N5�ܱ�  ��x��}���U~�.�s��KUaZ�y)������{��z�����,� Wt��Y�/��i�����l�
u��:�)C��ߌ�=n��S��y��u�ʹ�)�7��)��ݐ�*:���@�A�*�R�;�� �����UJ*/�n�$T�U�8�*?����4�f������<��~��
����M�s��O��3��u�|���U��º���G��8��oH�����5�VE����!�ns��,~��q��#�����[����#�X�[n���O�2��FєY�p�%�"z
��G�Jj�E݈u%A	��g�H7`ϭ�Za��*�g�[�!�I�~�NQ�nVh��ϟB���oȉsE��j�k�n����1�͎"�h)���J-֬St������c�mC.��}��&;#�0PhJ2c��<�O��VUouMt=��O?K��h��/��d�_d��Ja|_%p������ho�IÅ����b�@?�܃���2_f3́0E4��7E���}H$F�(Y�F+�U��B�&r6��I(I�'�x�B=�h�Z������A�IS$������,��0D~���p��ʺ`����*��|.	S��]I���f�a"���M��[��-��֦�*��k�Г�����=_AZ*�����Q��`�)7��V�Ô�q����I�GW��]6q�m�ь����蘮7[qZ�]��zrG�[^�h��ȍ��TR/�x祇��:w��ٽQ��� �X콙|>���G�֜��������l��=�j���0�t�E����ٵ��w**a�+Ӕ�ˡI%5�[J�j��%�e�O���]]�5�K�3$�w�ޥ�����c��>ߪ�ދO�V!m��fW^9�|H-�U�`�0�6�arz}�G6�娶CŇ��q�A�g�R���y�Ҟ4���c���� ������SU=t��To1�%H�	�V�AT�U��Q�:C�)l�A��K������+q�B�.o�A����'bZ!��0*f���jB�=ULp��㬗��jM�b��Ęq����R����,D뼛z�\���>x�K&C7�M��L��0�p��lQ�+�4�a�,:�,s��)�|�4y��v�� ���'�p@��N�8�f�n�i#�K� �]+ycv�UBC�m��qi���UL���c�&\h�z-:���y�V�������ısx��I�@�-"Wm�Sgp2�y���Cm3�O��������
���Q��`.D���t!��A���VV�'�Ra�v���n#�[����
��9\��p���r7��x
��	�6�+a���|2t?�P�r�7�{tR�We�%o;*����K��9^I�����8,Ax]W�eBO0p�g�����t}ȅ�~`���6��-�`i�2��g�B
��h;�p���wty)��İ5e�[���z{�R2P�:v.n}EVs��R �'���N�O�m�z"*Vn��h�Ӷ�T&6~q8����.�WbNV��v�ubň�e"����L��>�^��ٙ��:��s������m���_��)���)H�kRj|ʞT��ݫ�)8i�� y�Bw��o\�˅�R���s�7�@�����0��iF�?��l]�7���|w�����+���@��$����4�R�Xם�XlRq2>�
H�Z��(�^ڰ�ʷ�_�N���x��tT�G��EI
���˖���,^2tI�ƅY	�+AM�[���j�DN_|�.������>�10
���@��y�y#��Ks������F\�y���Wl�?�X7"�'�Le	Ie`������Z@��XlxVHYEB    231a     6f0��[c��Ȭb<Qɢ�E��@�O�|�z�q
��+-�֟/<.��4���i��-F�XCl/?����0ߞ���zqj#A�[<�[�
����0�sO�>?����q��7k��*��.���.sj�g(Gg�{��FW��꾁�"�J��0�*�nOd0��������'#��Q���J�$����I�Q�s}������������c����jq�7��X�B�RiUA��ɐ���J���AF���+a@������(oxM��N#�׃υ�KdB�����^�ԁ� 8흣�6o�U��p�9����i��/U)kń����3����m��-�!<0���gr�/~�Ϗ�u=6��H't��|���Q㔱��		՗9EH6_�d�Q,�i�J�w���&�qE�?I!�U����˫����h�4�i,�s��# ��΄f���VE�6�Iu�[�`k�ۗ�i�V�+��Mj!h���H�D��s��厩�QY��p����N}s?�Т}����ga� y1�V�g �:98��}�)��.I�b�Mo�=(l_\�h�q���i��zT���!)Зc5�`Md�A�(^�&��m�e!���)�B4Fۿ���Ύ?�qD��n��ę���@�{F0��Zf�]��P^���)2P��Y�v���7�k�oT�_�y��ׇ��;����T��+T��+���@�|���&�C}T|�&[�*锐�x���/w�s�2FE���$*�M]�7,F��}��bhg���?kS "�/?:���4�ţݗ�#�$�Z'��&�#>�Z�C��j˛D��9J<nM�E�Q��q��F��>�z��a'�h~�+a�B��I���1��\ &�A�A�'�,0Q�?�6Q��/�7þ�3����Q�C'�|��|Xi/7]���"*œ�;�xKz���_D$�<�d�a��2��}a%�o������!qҎ�1���"92���7��P�����?b/N�QB@�n@�^��D��2�}%�LQ�[�Ȳ�7˽"�G�3�bb�����*6Jrݡ�Ch&��k��l�S�/����ݫ~��L��,�!�wyi��j8�z!m�4`G��;��]fkP�����K8�y�uvf�r�7�`����s�0������_-�<�Mw�i�~�`�O�kM�.����l�ՙ�Ɵn������<&��(rkIĒ�>�Y�wm;��b��+�C�'
[�(��O�pF%��Ҙ�Vp��K��;���j,�'-�R�l�<��iO����A�oY�}N�x9��F
#��P�N�~��گL���D�NO�֦�-��!�e��g	` �D�[�5�����v;�~�F�8;�\�n
��Kwpߓ_k��/�寳���I�9i��ֻ*�Q���.�����N�t���H���]�&k��L:q0o�1�b��caF�SA2t��Nw����sk�"�4���}��шW� �~@��
{�	K�� ��Q;�S�)T�.ߜ�jI.~�ƿd�V0 �eٹ�X	���@���˧�)�Y.����76��)�,��Nb{�T���T�_�AF��e�c}Y]�9k6�%)��L�������3{��JT`�tu�#%�����L�^��%|�80�@f��x,b�1����B��q]K���I��Z\���KO���{��>�b7�ǩ�A�xQKi�zҟta���ueӥ����$B