XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��B��ss�t���ݤ6��Z���]�IYEs>}��V������#�#��ds,��gx^�a$���H��N���δA$�6�P�����ټh�u؃#�O�J���~�Pe3�O���[��<t�:
���G���+"�Zq�<bhY�M/��� \F��v5�ya���Q�i���������(YŽ�Q����DYbo��	�R	��*Te�o%"����?�BWy�U�Dh��<�0H�i��J��҇��;��b#Z�'��o�h����JbbF$���6ڈ����1�Ӳy�h:� �i�eÁ{΀"P��,�2��Vܥ �p�ME��<��p�(�
Mm����8��8o
�{������>,ɠ$v��7��~�M�i�|�ӌ[*pY`����[?�nM��`M�"߰�mMF��}��1ˬ�)��3���xPIs�`, ��
#/me1v������Z���w���S/�̒�Ze�1B�C?n~�9�����j�SR&��s�(�E�ݱ� C��fn3��[lN��+���E��O�oz�[���UȐ;�#[�^��|wO*�R��LG�(��鐦#�IR��O�ڲ�Q$b�_sU�,߶��!���gWY�2<�K����Qb���D�r�2B��d"M��ᾐDz�g�<%���mt���#l���ԯՕ]�/V���I��Y�~`��0WeGŬ�;�� ʿ��FIf���_�MC��`�և`*wf5k��&��$e�'��u̇��++kXlxVHYEB    fa00    2a40:g���I��5�� �#�a�����EtiĒwtf'q-6�uv���:�M
v�8��-J�c!��c����w� �CaXj*{�V�%���J7���Թ5oU�u3魘�\k�h�W.Y�z���GY~�T�ҋ��oǑm>���g�����8�Cغ'x���%���i�8�ܡ��dz��f�'�~���#U�N�ȁ�XY+I!M��R{Z��:�@�+,���B����h �T�'!'��"E}��'�smM(�h\~�9` ��pw��6**������aRB|����I������`�[�\�h�	�"��:n�=�F��'2( �B�W|�;�*
��-f��yD۶;E���n�iP�z�ل�8=27���w��-`���dyb���(b�ɏ�9enVC� УMu�$n͛�jf�q��U��k���+�<����9ɕ>^1+l�{�/F�w`1�o}�Z'o���/ݠ��5�*�X_��{�WQOδ=9�Pu��`)?����v�� �
���{������[I&~xYo6�%��!E��b��L5�o��,�cZ�����A�����٩�^��X%Ë+�+c��\�~LJv^�!��e�#9"!NJ�q8~�#�*ւ.���|�*]?ݫ+�T��$!Ħ�53�H���H��n�}'�ǖ���ca��im_TGw�,�;4Z�	��QI�����H�h�~)�#.�]����C���c2դ3�\Ab'��o� �),�-D��wv��H��,�k ��?Y��0H��.�w���S���z������C�8$�6�ۙ���h�@�|{��7���"{�������j���ۃ��M�������"�CP*�,��ѯ���e��+�\�D��p�=J%��#]�,�-m�Tf��+x���J�-�����dH��`g�}G@�Y>�H�4��Mf�� t������ͨ�Ԇ��X@"�~��E��Q�
��)�J�e��l|3�b����~^����En0R��Rj+{Υ���a�>ڮWr�INU�3qEİ�M9�_��2�B��`{�+���Ù���)#go�%��Eg6#i�Jq��=:n�|��F%l��k�.�%8�Ԉ�}x�Z.��e*��:�S�?D�7jU�ǮXӼ@߬B��z�U;���.&-G�e.���n��E��
hqvy(�@�k�8�,>�_Sc��b�����U�d ��� r�z����)�`�\EPJh�:�p2��cꈪ\0�4���/�j��� >��S;W�6h�+�K�l�.�<��#1!��=�M���T��`x?Z%�]ؗ��P��t�O0�3������)�a��5 �3�����_B��BԲ����F(� ۋ|+���]�9��.�5͈�|AJ�fִɬ�}�z��-��x�e����)���� C<lV�Rg�,`��B�w�wg@x�o�H�B�C�����8"Y,�Q38�8Q��N�N�-�Q�Mkd��~ݻח��38����Y6��|Qp�wľkJ����̻�O���Pf��'c�(lQ๎ߚ��n�6��޹���}?]^����m�����,��F9���ǝ8�t%��.�<x��0�{ �c��dTc�$�gW�M+�J��w"�D�˜��rD��7�m¹��W��;��'�j�, �drc9s{�mc����8<�5�0���L�]�!CQx�\�j"
�;�<X?�VDIc+�'�5���g⠮R��툽�/���_$����En��-w���jbHjp۬be.5<��bt9��U�,�oS�:��r��FK��t��Y��2��(d��Lɲ&a�I�XK�l���EWko8�m��t+ֿ�R���a	�Q��1FO�FT�:���~�����O�*o�=^�&���Bs�]��5K
�:}�>��O@WP�t�G���M����q�1�E��Ҳ���>"�@���H�	C�@�CL���$��,Ql{��g����&k�5�q�`<H[��]vR�� L�7T�P�}��V���T��2]2Buܜ6���~�l熾hj�ўǱ��]AH{��^I���c��|^� 2�O���D
נC�>��b��i|v/�$(#��%�v�Z���b�����r�:9����);�#5��=6j��o�l��!	��>�V���wɜ���y
"��<F�wu�E��e��m�v+A75Ϩ����)�=��S���{��
�yM�������|󵎠	�,���@U������O.W=�����t�ϸ\�q�����1��]'�`Sj��󵓿gfݽ�k��=�	�V�jT����I�QByp���[c��w� ���}v]�)��kҟ�&�l��4�AN�5F+0H�C�8��Pұ����:{�ܒ��a5uF�>�_����Ôb���v�'�8�=]N		Pvg��x3��dF�V^�购�[���@
�(�H�548�����H���4�s[n*�R�C&�
�v��������<i{�.%��nq�9e�P	�)�*�����QNp�H�}���ѥ�Cz>>o��l�wC%��T���#�����mN�FZ��)��S��|xGN��S�������
��Y=p��HĞ� �&�@��E��(Х�N���-�i��X��4	�"ۭW?E�<H�#S��E�T�צ�E���;o�+�z%Ơ��j&�l�@�1@ِ���3_�}"�tX��/S8�5�?��X������������Ng]mō*�����G�>��Iy�-E-�|�b ���Q�����GT=0����f�r�ޑyueF:��k��I$E��40��3S�#�Ǿq��T�X�����/�9��32+:qi�r<���=fS�-����F��܇0��pP��/pz���[A�A�����,�O�7?���+k]�=��	�҈<��ɪ����-�y	c:�&S��J/&�}��j�6�C
��'���pY�Pɛ�R_I-����;ұ{� �B(�h:��y�]����z��q*]���/�4c�pcj���N<\��?��LZ���iI��`��h&���F�5�&�<P���?��9?��agB��~Y$�m9��SDr'<��1k[��<�����Dؿ.�c]�
<%}<e��F�<�*mY�X7
?�iI2�U��oQ�ݾ����L���㥱˛�X����\րH���l�,x2=>���$NQ�����q�0bT���c���S��Di���
����kh%��Xp�-����V|��l"E�����&�@v����`J���F����n���6���������;��M�84(��6�B�
>ݲ�l�k�ڇ���c*,<���4�nc�F�� -��+2�Jy�P�m�%f�H�a���*�5�dt�B�k�Ӵ��H�`��*ت
^t��+����( �޼�yK�n���a�nii�Z��ȇ<}�\��>EM_��		���I�QW���cկ��At8�0P���/S�?�z}�8�[c�_d铂0EP�oc��6�d����R������کm���9q�3�=9K�c{XP<���V����UB{CgΨ&ʛ�e=bt���F&%�r��
�.A��_����#�\�Ƙy��|n�[
E5�[[�Z9�UE�7��M��O=����N�3Cw}76g ��F��ӆ��S�1{z+QG�����i��ou*��uHZmH�}��3�8ic%;�:���g�:�]MyIt	���%	�j�V�Óp��+ ��.������w�E/�'�4���^�j�V~�H��v��Q�~�ߠ�v�PދN=eW�ܶk�o�&DI�n�� ��D�!��n�2J+�tH�_��ZzУ�[�J̋��"���{��l��f��zY��x�yI���i�����=V,��/Ȟ��
��F��������J��`$D���'[������D0�6 2���1'��O06�9��V7��D��Z������`^�3{X�V�=�y���'���!
�#�;X�y?ǖ8��?��������Q�J�S�-*�w,�����U�jj�R`4��7�u:N�y�hN�
��0���(�U}	�ꎛi�����P��b��˘(� Y���]w�C�����Y��\]�!�b��%6��I���/��rT�
��R	K��c��w����a{|,c�9���m���3 ��HZ֟q�F��_��3]��{C[�H6���Y&���l ��~��,U"IKS�I<��ʡ�߭ݱ��������x<bz�����+g�5nr��?��%���.�E��	/�cIk95�K9��D����Knϯ����mi���+�]���X����P�GWS{J)h�F �C�e�Q�C�
{h2��T�u����;�$�<�fS�T�O��fľ?����EH6@:p�s.'�)�)�����{p8ٸ`J���P[
	��Y�=�����ӛ�/Xg۾����F��k���d�G�b��<E�@�T��Ė_����k����^�W�u"�22�n�>���y�<yS��nŌ����~?V+	f],�n�DC�lk�rC�xE�ewDk/��R����a�=3�rM����M�|��5�)~`� P�_�������j�t	Mn
��s�c4��-Y��ک�(�_�����lO"&�5�A��G2�����ML�������mE$T�e�x�~�N>tݨ�?pn.��x�lZ@)xN��PV�0�O󙮟�qi#jV�%� �͔�Ж�?ZI��ܘ��,M���D�l�=�´"���H�sQ��> �W�V�TkY-��آK��V��T�n���ӟ�}k�s8���w^I�EW��g��{�^&]����/#�u/j\�G���A'u�q������	���Ïc���dbѕ�@�`�'Zuψ��
b��	�ɩ��b�E�3�&>[���tY�R�F1Ӧ����2es1%ѹmY�6�]�/��U�#59��nm�M.�"D�h��Kv������� sp�ɓc8��˻��v�Ҁw�Ψ��Aj-¹i�}xO��O]}�F�(��3 ��/��59b�����M���C�M>(	�D�_KQ$N� 	��m]����jp��V��;�v)��G�Wf�K���(��<bS̒t�蛚t�nظYl���d�65;b�JSn���˕ڏA-����](�z!�����B2�.�|�	M�Z�@��觅�CD5�O�o&���p��\)m�ex�~�u�ʨ��sǃ�|�vgo0�`�#!����$�:����@�\O���6aP�} ��nPN]i1�
+P�5�aKZ%�I�}=P�
�{�s�r��f$9�u�oľ���,�e<l�7	6�v��jZ�Qs.����Y��R�Ԡ+��O���ኦ:��gB�y>}�xVu*hE��7�k��k��<z����EY�ӧ��4XͲ7�M�jQLG,r���>���k.(IQ�Al[�g���*�a�N�i8�
�����t{|�CvK�8K����yN�c�3e��64���7��9W�,�N�[)*%)��;!���+}�T�J��4H/fo,I#����Ը���e0k�$�l��']ޙ7�M��S<!]cf��m	�V�	�m�n|�#�:c_�'�ms��8�|#���N[�c!
#��8�&��Y��7#lok�\��((�@bFZ��,�����4,�܂�$ |��:���t���w4*��O�h����c�`-�v�����ޚ�Xv��D="E����g ��"<��s�b�@F�+ʹĉ�Ǣ���ry�B��toԅ`��M)6i1q:S��dj[%F��� )0�,��]�M� E����w�c��X=	�w1X�[D���u������\�����EY���tMpR���L�[mTJ���c�6���Q]咚{5e|}���q1�D�l*O�Kr{�RZ������ �6Z,�m�n���C�w�7Џ	l�a���S�A<���4�����F�r��I
n��I�j`�"�Zv�V����R?��f���,�&(�jyDS5[�1��8�^��^ݯ4ʆM�`����
� [�y��.��m{G���׉u7m)X�M��� 	�z�&k�>�.gqy\a�l	B�`�� ��Y*�Ԕɶi�)���.�X翉0x�M5��8�+y���r�IC���w���M����*��s.u_ ���'c3E���o%"B"�Aܐ�ִ��1��W�
s�d��ק�����㔴�V;������~ l6�,.�L#�q��&l�����@�"��rkp��&п�0��5x�VĽMe��=q��˦fx�����G��7���4��(���*ye��7��5�a��uC��kw�k��fR���0D^a �j�X���.=P��x�ˢnݤ2jxe�P$w�[ǰ8׬����9��^id���h�^ɰ�6����֖������v�F������R�)"F}�V8��P.��,Cϸ��_�K��<r~�kͮ�%����m�w���SҔP9�oɌ�5o�\\��k��5��������|9J:�C#��ʖ���ky$�p�.�KU-���c��%~�
�FC�|ޥ^?�T��#���V���;Vh�c�z+?��S	:~�^~���!9�$�^��~��BoS�\���h��n�o�����f��mI�����05'�E[{�����E���7tN����DJ���Ap��B:g�pP�m`���L���yd3r=�K~F�<����P3���1����+ihDJ�ŽW��2�C��V�?,����w^5��-����&��gsR����R�g6��{��>$���ę�l(���Z	����<?)�Btenj�iY�8!�>/�ō��;��l��^�[�[ЎRX$�h�i�5���.��7P�<&zzV���Z�T��&D<���};l�����D#��ݨ�kԚ@�7LX���<ه���ڤv��\2z�HX�ݝS���Wv�>$^V��D��q��l�.����e���{�s��ے�t[[.��쫎��"2��N�h�#j���в��w��~ �Q�G�]Ӥ����"l0)�}����?y_YBU%A���!�LU��.`�/D�d{I"0%���x��wX:�3����'�K6��Ki���mK��1���Y������ڼ����a�g�Mq�ת�N�3�b���,.7��y>x&vЕ��F\(嗮���c���F����[���dW�F2^��8��� �q p8K+�DX�X���;N��j����U��t���o��&7�B)O�ᖒ7�}����(��j��iJ,-O��?I?p�9�@}�[gɏf���M��MP��mx/���򷚙��G}�4��8R.�7������G�f=�/�7����Ac��O޸�xo>��fTi�yf���Q~AP����o�FQ~�</{M��H��m��0��%�]���I��=�!ں}� {��$��o��r�K*H��ۇp`T�Y5J�	���­�Q�����e�8�T�
[
�����ŧ�=�5�~�X��Ul
kU��˥s��T�*�_B�r�Gm�/v����@^��#��<N�����!u��"�����K�)�/dxw.^���kq׽��Qi�W��l��p��Q�W>_����/z��6<�����!�I<�|or��J/-"�!������O���(;�9��S�{ q���Ӿ%����/-ȿg�aw���w��>��}Dr6�".0pU�`|U�'�`��"�.��_QA�M�?d)���B}�֏`��"��х�yD{0�o�R��@���6���
�;|��뒭��\�*�bX�=��%�����R�/���`��}�o���W
�J^#�r�;�-�gK���X���̽,D���>@���|P���s3�wù��;) q� ��8�1���y��h�V4��x��Z®('�?���YB���6�htQ�?v'/Ugհ�Ys����j�G"��d�v�!��F.��O�G�p�͋����y��F�� <-p���
*]�)A����70��#���/�2G��߂O��RF�d[�2��u�2k��(_�����$n���M�9/ӹ�$��� `�>��<��G�Uz$$�W�O'� n+k4��5^��6Z�eP�Deb��8:��]�'�;����Cz�:Z��ӹ$�hQ`�������Z�	��fvS#�����ݪCV�X�������&V* c��\`��1���k��.�k�:��E���*nQ\w�Ӭ�վ����!̛�g�'P���؎��[�ݐ�ۻ7�<��}[j%8b)�y�%�e�o$fe�=f�T��ms�?s�G�
�/�>��rN��H�H��9ac��G?���S�jn���p���'������.կAGO�I�1v���|XP2x��TCLyd���yn���H���V�W�l\ű7SlCkً�28Kj�Ǽ�O����Ⱥ�#A��%��"���ad�o�W��]1�x�$Y"���/��4&4]�����r1���v�l�hsCf�~��o�K^R�/��.�gr�����=�|If��_����5��m>�����+^��W�x�n���5t��՗�Jdq��K�����O���LHc-Ӟ��M�o\�;��>��&?݃�:I�CD��ʝa�xɉ:Jo�#�bo�>��8�"<����{��;Z�������k,�B���M��;�w�:`��*�2�@ݸ�*���5Y|Pw��V��M����� �9����h���2��|n�A��$�����������Bp��-V[)�x����u�Sx?���@��z4]�(��o,��-7��+M8e�K�,5��s'�2��٣���-~��co������t^g�����p&���U�קz����G5>W+���T�2�M�o�M�[?��16k�S�V%��Ql��<��qFdr>f�)��Ew.�I8�@)q��?��En`?�M�I�bK�DFr\���� 66Ŏ���[�=��=àSx�
�ʹ ���"�C�u�io8��a�0�Xi�TLS#[��\��v�1�R������Ԧ�š# <:����{kW���1��×�~���8�Z�ґ@��}K�7�5k��	��� ���_���6��p���;ߑ����z��~%�ЊO��ځZ�/�T1|��g{Y�B�N{.5Dr�;c2�fvF��c:of'�[�q��rR@�T��M#��6��-6��Ȳ��3�G�L$Z8�i[�����^86��/�X��]J�O�o�W,�V�ڡd���@�/D�d� ��l����%��g#O���W���A�?��]�S�b��0� ����_�?���,�(�_֠A�4�V����$�a�,f�}	��Ro:k���O���ہ��B:�ҽgw@��G����l�;��n�;��D�
\���������xv{���`���bL'B�j�r�|�ޠ��Ǭ�Sp�YA�;�k/��ʹ�F�!'���h�ތ�2���Ys?7Q��Ĝ�;�Y�!�4eQL��`
���+j�M�NB���{�����ph�O����d.�M��)<�X�B2Z�T�o�f»l71���H�Ӣ��X_{�m�ce�띿��F�2~�`�xLoo2[�@P�!\>�L��NM�L1X(�Y�"�i>�f�3��Ɯ�`l�»RC%��Z+�Bd)/�3�.~�ee飫/���Sb���"buL���v=#�U���3��tq���\0�?Q��w��@��e�#�՟�m�cU��ݾM�}����N�(0��Dl.o�G�����K��jR�rSZ�t7(�Y�|�KJ ?d���yө=�۪+��9'�n?=#���gs�1���Q�|�ׄ���6GZ�C7�`�~'��q��xz$|�6�mb^&`xVˤ��Ǯs3NC�(����."�s�o���)knf�|���:��o�P"O?#�w�E��]`��&�<�A�QfJ��&��`8�g�_��3�M��8�N����ʇ��$�75�R,؄�Jˀ؆#h������0���k2ކ<L��K�`2� ��e���=�t�����/W��f�G�{�1hu1�vb��188Pz�Ap����^��#=8�]��>d���R}�`�E��G���j5��fګ�g���ak�Ϛ��wg�QV��^�vI���#{�ߘ^z�E"��fQ�Ӫ�Eh6�{����x�P_*�����R�Q�h"�>�U��Z���Dn����x������Bu�mbk�NS+�,@�iTLL��'��BT�v����h���[2GĄƼ�����R캒[(h�jL:\�������?�ͮ�p��v���9p>ޥ�u��	����NNG�z�'��׻t�H�ͯP�03r�&�%FY���j����a���Fv@�1�\%�5+��ϊBB��Z^�ג�K��9��M���;�U�%1�M��0L�vm>w�Ah�a2��������N}��}!��E�̓�T����q�H�#�.(��W��2���:�+9����2��y ����[��Qơ�s~vf�4��g�#�r o_�����i�S�4k�ӧ$�*!VsI�Ŗ�h�
��:��~�[&����Y�]�{[�ZM������w�s�XlxVHYEB    fa00     8e0C^:���ۄ ��Nc�����x�>]XޅC��H'ckTu��B�F�D�?9��H<�i��-��S,O\���r��ې�.�-�������]�q��dAw�pa��z�7bՄt㙿f�6/g��� �$���7�T��7K�;c��㬋B���^�gL��fk:��QvJ�7�@6���ln3�������{��������t�������e�O���x������a���t���Ac����1V�A5m=�Z�H��u�ձ���[��Cb/O�z(Uч%�3��r�rKw|�*�Ƽ/T�����*o��5�'�i*H�et�ŘNk�1%'�'���s��<3�Ԥ,	����03pF���-A�C�l�Ge�H^���L&�*��
�$S��7P��M+Z��_䦨��P�l�痌��A�UI>mX�x�\3EhnJc
_0�"f�a��эw�Z��1֍!q���Ar�PYؒDo��z�y����}_�U��l��{�D�Ɂ����~z.�,�)�Ɂ��0j��qR�.3K!f�c�g�am������8ض�k��Gށ��ݽ�zW���I��,�5�#Ya߮��,Z߭17'�z�����*���:���-Y��R%�/�	lK�k4��P���z���|��%7x���������wĐ�j�4RMդXUkC�"��P����7gu�K�=��P�%\��?����y%jRSR.M�j��P�j�Є�#W^�n��O.� �����[�o3��v�H2#E ����vZQ���q�S�f'w��u���%�U��{�]{א�׆|E~���gf����ݰ;��ק��b Y#k���]��4� �|"{��u���X���Z�����zĂ���E i!e������ ����@E�<o�L��P�6��"��c��J}����tі'��*��* ?�L��k��`�b0R�e�m��b��Di:�ev�x�9�nA�3"�\xS?7~9}������k�6�Shr6��*f�*��ֶ����#cV��3��Eb���_���Q6!�9�d�&�N��g�S�w�Y�,�]��^�:EzY��+C_?zf_�$��i��hp��MA�����^�Xh�DOV�Fi���������!��Ms������H4}t���x����K����f"w���%rs�hBhx�#}��_�-mt:��qO$��*�0rDv����2��AC�}bL73	�L�y�t���'v�c򅌸�5�Ռxe ���؈�]�Z�5�:��hg���0�f��G�vr<�"�����a~yO�퇁W�4�b�,�+7�*��A��j�n���7Oi��ɞҶ|o�\^It���~Y�	�
�\���Pf�*/�ŉ���'���0��4`��0�>���8�zf?�W��l�VT���6l�R��z�87l����W�͎r�~
�+�F.ƨ<�x�{�&�2��V}�G�#%M|�wJI����r-LX�M9�bh<��^��=(���|��s7�c�c��º� t��V%�L��+��n��N��E�����<��דT�>ᢾ�g1?�;��%U��W�%y��~��^�$#�	����ͺ4w�	��Z2��"y�j�"��s�V��J���Q�5x0�.�;�_�OV�$�Q}��	�J��	�Q��N[����p�eR�,kכ��K ���*�J�E=��`��9D[��wd�w��z��k�Ʌ�rD/K�X��ާ �ɀ�w�T2�Z��L��#���C!0x��ޜ{���N$Y��	-U(�l�'��+T����. g��%�~����'$ث�<Ѵ^(�'��v��B��&�o�.�ªօK��扐�I���י�\A
*���#��>�9��%��g��q��4{�oa2��lZqb���|k��O7�E9;t��)��]�l]׸�~P͜�cI�'����hUX��{"'gX�S>���6�-�:�
������a&�b��B������q,�6�Ħ��>#b���j�<f�W��������%C�/�'�*��	���wl�ݠ��Q�	�	,[�'c=��\�F��
�X�^�0���o�+BF� ]���:���7
A��b�Cv��u������?D'lg�D����3�HP����L-wv��h5��3�ٿ�
���"E�5�*����9��ae�B���Ъ�A��.%ͭ� ����|"\"E9� w@��<t���[����[��^\d.@K(�ժ)JH)gXlxVHYEB    fa00    1110/e��%|]�!��(��ۮ���Vƣ'S�5�Q��5#�����eV���RV7|�
��t�HH�H���O��X�V�K��2޽>��r�4`�d}��d	#d�Zg"9>X�J�i����J�\�,%�*+3��lUc����x�V�qN�1(#6���I�Ln��	��;�&�m`]e��Q�U�@a�	Y6���6���qB�v>@f�o�)UG��wDDg����`��3��`�Ji��NeP[3�mh�_���	��m�<���f��3�(�S��wߊ�(M�ܺh}]�J��D�+mS/_؟�Ķ�L�EVC��(�M#����7��e���n�6L��K�Z���j�뗓o�� ´�j��PQY��c�	*&!E���B姀q�<��D8���R�:���)ݭ���?��n���eͨiT��ٽ�*���3G>ȜE`Jt7<7qg)��l(���i��3�����������(4ZXsK��ӂ��+٫H�r��W��p�~�G#�������y�R=�r"����s��!��N5X,䏺�wgxp�əɘ�����%d��`��X����������"}����l ��ɎJ��vf���߇?_4SМ~V������R���k����4ѷC�H��|��4{L��T�Z��{zXwK<�7������`�6�Tۭ���Dz�� WZ�Lq���]�u���2�<
�f]��w8�!��w�Uq���b�k�RGA��Y�9:��Z�̈́y��D+������2;p�5��	Z(���T"�iuxZCCE:J��n���&s��iC�����9�:Q�T(Y�B���/��X�J��;�qf0�pǗ�]j�R
�p�8c��<4�{�
���&�tۨ<�>���%���
,9�XK�����`�ص�[�[����= ~: ~Q�h\�c�`������+c��^�\VS�����	������+E�p^��S�BB�쟸kJ�*����!7M��W.��T
��	�K���[�o`�'�wc�J�2�{祔��w�0j��s����ݪD�hw�/�{�� {�"0S��L4���������ɾ�4x�JP.*p�)bl�.X�]n;�Y� ]�9�a%p�Z�zb��y�C,8�h�q�.yj�ЌAٙ�^A����>~V��={�*���棏8eu��Y��$nh��_���M�nY������/k��Q_���ؙ�
̢�cE��暶��~CIq���˱?�v��(#�;�uf&zDj����(}���)"��%n�:�򞔍m��v�`���k�� mB��N��( N����;O�#hL����*%�3�?wh�0�կ����vRs2��kU"L�RH�~Q�B�iz^��5V#�-OR1���6W�C��7U�+����"2�'ņ���Hf��Όй���
��'��S�)�����'_�Ȓ�����Ny�����L[��"��v�,1���*�Ԭsc�/on�ǻ�`E��e���E��4X���rG��W+UM�9K �L|/���v[�M8Hh��Y��fA����nk�!;�a3̢�Z��8WE ��]��y
�HM�IOw�U#</+��Lv�3��x��� r�K���#&_�v�O�q9fW5�q9�=T�@�|�� 5M]a(�eȀ�p�iC6�ĭ*jL=A�{=���������g�܄a�?[�=E,���=��M�kQu(˲=?�W���]i�M�i5�L8����l�߱�L/F�C�XB_jvv�L�*>-H��5PԺd3��5j��z\��p+���e���n��,��������|	��g�aDe��@|�'�KN�&��k�;'4j!3���?���b�����b�^+�
��.A�]��Cnym,K9Y`�^1��*@�+șd����wQ*�i؀�Z��Xko�����A����f������w���2a^�|]/�+�
X�Rf#B��pav��^�~\͚��n�6h���	E�0+^�QV��4��*�X�����^��0.x��A��.��`?�~��&
覒*'�ݭkA�W%��ix�\仾}AD��E���g��p�g����Saܕ=��,�;�9�q/"	�cf��*�����E�c�ڧ
r�� ���U� &��b����D��b�Tu����i�]�W��w�c��ƽ,���M*Sp{��I�����E��'[9gL''�%ڪA��yؑ���Yr=^.(�Z)'�՜�>�<3�O�-�T�L0]	z2>PhԢQt)��>�r�;�?��ɾ=c落k��ԯ3���2�'w���ǙYs������
b��ں{:�R���e¡�Eq�	_��N�7_B�T�!Cp�F�����NzGW]�=(u���\fe���r[�H/�T�r�!$E�0������$�
����l5F���&L�,,:�Lق�(�p�Q-����LW���N�t>�CԐZ�s"�H³II�yӑqp	�Z���f[�ǜ3�@�ˢj�`F#�Ῥ��J�>���bq%ԍ�>8���p�/I��x�l�R2����E�Rx����BA@o�՝?��T��&�e�:�|ViftE(ә���/��9����P�����&Ha�hU��E�(D�2v��X>>{���T�� ��%���i�+F5HY�C 4���7��N���C��a;^�=v���1�4��<�?,�w�Ѓ�!�#����D�T���
@V�o�h���2���XI��\M���R�q0CD`�/>�`��:��Q3糆��L��E�*��)b9��`r;�`�u��q�]r��q#�_��)!ظ��"v���W�\��F����bŇ�3�+c���N*$�Wp�mQ7�I�������7�L(�~e�D�+��ӆ�chYF��5�U�΂z������3N��R��s�m[wFc�E�7��֓�Ӊ͎\K�JwO�s�ֳ��`��b��5]���3���6�j�n'�8��pn�,=�[z5ق��ׇC��f5L<7��r�h�=֎��c��td^W���ENj�Lm犖�
T���u�Y�olp0�Եy�ֽ7`���`<3�!���*mp����.|�f7=�3��9��j�)��}���5\�Y-T[wC�7}^�_�h���@%6�9C�Sk����r�ٗ�,���rX_��g�]ͪ��?� c]�B��	���i�}	�Z��gtB�`��a�����lD1F������2��E����� ��z�#َ�H�9�HcO?�y�h��(I��ܰ���N�b'��!��w/i��JW�m�f�����3"�u'�'~�0��8���]�`?�dy���GG5�nS|yJ	�Q�7z��Ӗ��w�s���t{Y^��3�>�I}���#0Ȅ �0Ϭ<,��mq�c7"`��*4%��qB5�����U���5���3�beo�,�����Mg���eI7:l.�_Ɨ()=}^�g�ɉUJsa�w�m��|#8��/9hJ���GPa�W�|lc��AV>�d�����1|t����ƈ�>O�O��X�r�f����`���_�z��p�F�Ib=�(ɔKCs��ĩ�����N�)��y� $ �N���Ѝ��/�G3sm�I��F�4�j��1(E�l��I��
�)��K�3>z������w��� ���<
�W��<�MY����W0��,q���h�����y.A����y���ei�o� G���uo ���&[@=Q_�Ԥe���F�Tʩ�ͨ�P�~#�>�B���)��i�{m^�,��CD���7�0M���b�g�f�|Q�~�����|�l�b>�����%��s��g����SW���n�t򙍵2��d�Ԕb��5KR�s���B��|"*�?�#ֺ��1·�Nv\A�u�t��5tX���l��J3��P�����q��7� ��l��&�Lm���S�ۡ&�� OZ
���rKsB{�t�࡟J�	����)RP���p}J�,�� D
��v��n������yLm�P;e�1M-@����^hBZ�UDt+���V��)��a��y�;5|(&�OB@V�����L��n�y.'�\�]��{�R�tM51��=�!��?����%�xlr���`�OM4�RyR��Z��q��Ǚ.AnAo#�Z^�N���G�UpPm�sY���<��ǣsnć���pU�N�k���a�*�N�	wԝ*�bAOk�Y�O����]K
�����GN��y���J��!w���u����Q�BhCR�.E>�.4FLB��+��aݻ@v|��X���XlxVHYEB    fa00     ca0|�¸�}7�{S�����{�.��Rop�����o�"���y��`�bdAL� |z�iY�d$#�j��#*آBQ�6�9�:;����ih p�a����bJ^r���#]1qÙ�lT�vo�Sķ��0x8J��PFJ>�{5I�s���8]s����.��@փ�� <M�U����|��0�c@6��T�q��d8ύ�x��7F�R�:c�q�X1��n�;��
����V�x��REY�v�%8n!�4k�����mAwz`V�<N�������y&���[�$\i�f��C�L�	GU�g���8������xY�(�8�*��dfИ��Rs�'ZXeu#�l?���3�}^-IJ�`�=-r�Щ��gF��xy��.��.J���j�^٣�KG����
�
Y��FvB�K�:9�S� P�ǰ�쳒4/��Z`Ў7�H/�����#sB�-r�BWg���M�b>)�^��S�/>�ޯ�+�dZ+B�>PT�N�Rm�Y����þ���[EJ%�rJõ�ӷ�ʃ"������+�!,���@���ȫ�:��P���t_#j�g|�񪻞7Y䦷,E��4���	��+K,6ˌs+�w�@�w�Z�pG<��8� ��L�]Z+Hw���ZD�g���]�)ӏΆ`|�^Lch?"E���=��vA5*'�m:奄���^��V�T,�d��l�b�׽�6���RLb�������U��j���kP����;�\ew�ǧ#ec��y�8��5o	�������i!O8�ߨ�D�% ǯ�Eh'�����["�]������`^�i��?wW�ph��-�������}���shIca	��\T�2��6N�H�o��:���������L%�b8|��2T�n���ʮw�s�p��%L�8ޓ�����=�̯��{Wy�Z��N��Bt�;����dy���N�Y���.��ݔt	�d �n^����K��8'�Ƭ|d��NBZ�p4����-�W�.�8����UR��m
6�[C����,@��G.c:Ri����9O�.�����	a�Vh%��89�o�^QȊ��ahzj�/��F�犬}�~-n-�3�꠫��(&F���g�Z�*:�(��~6��6�D�s�5� �Ds���O��tm1���`�L�WW�L�0Q=��E.��gA����a�X��s��ä��5.�Om�r�ԕb���n�����А�'��X,����`i�.�L����� w�G/��ڴ)����8�AϺ��`����ؤu�#|��`;(���n�9����'1�������7�:F�?�nZ�1��.�)��'C-ì�&���N.��C�[���`=���Y֢��|��80�9Lu�I���s�O�j�a�`ɖ�]�L�J$}����@��ǡ�qz��ջ4�1�_<O+��\\�8�Ƙ����۩�2'���I�S�GU��-�����%�'x�����H��<�X|�鼁�U�G��mv���;Ͻ&t�Ʊ���A0�J)	��yq#�p��J����	ȶ���B�O���TY7ut��+5�FPt�+�K��KB�� �\V\x�ռ�q���Ot%*��vB�v��ھü(�踈R�n�O��oz��	s�2�эU��4d�o�*6]B����l���5-�$r�n�M��Ħ���Ka�M��v2�� ���o�b�}��6>�sd:71�|�n?���}�_���䥹��?_���Y���NR/{��y���f,D/�4��}�*�;�־��zQ������&W /.�Cא_�xc�w�B�^���#�k����bVbl��~�	�}8~��$�T�+4$���X��XN�+�g'���IZ��8�t��S�[Lt�A��.7�%�U֜���`69���2Ob�����V/"wX�\��5-8�ПF:oR��W���t(��ܧ��x�9F�`;Kؚ��w~�^z?����r�c�t�.t�ň(��'8���wql�����J�Q������iH�l�� K�s��0xɝ�֐�[Ӗ��~ 6�0��R�_$�ȴ��T�Q3n+R8�ڮo�5҃Y7O?���N<�1�n�	��q��H�V!��F���Oԣ��-�< ���z��C(zVp�����I�^�?�%z���="��#����f�j�֋%�eY<H���̘�9�.�����N����ܝ�w�"�Z	�����)K Y�dKz�%QĄֻOʬ��F�jj� ރy[�ZT��,�=����v���(K�ȮQ�t@�>�JR(�v#-�8���¢�5�t+�*B����6%��:U���C��f���,���/ڊ���~�pi>��,�G]tS)��|#�N�;��Q��"��"ܱ)���t�%��]�x�"��{;����j�)ԋ����Puu�=>-#1F�ү��]f��
�*1ڦX���D�$�ON��{�C�����Q�^�p5�ϯ��+u�=L���:_��(���34($�e#��FC�Y�lbW�F�:�A9�v�)V5�DP�¤M5]�V��©�N���{B~M�,w)���ּ͠����4�ϥ��e%���F�!���=�h���c�r||�p��l���x���2rU-`�	�ߩ��K�����ϴ���{?���2#��������M��o'��y_(	w #\�~���l����Z�ט��IQ���j��&)O�� �l��b^�T�$&R�W/�W}D�k�V��1�ЪnsK~�.����F6D֊�Fv*rOڣ=��o�G���6y`r��ڌ<�5n�f�r�6�XNC�z�ts��D~���w`�}��:�?����e�ƓJ�@���`kwUiQ���*�+�����|z�%Ql8O<\Z�a�N��j_�cjjd��%o?q^$e����n�h��1NzQ�;��nrB�e\�=;lV�4��/�T��.r���Q1�gnh� ��H+�� �ao8������;ga,���:�����k|	k��� @�/��d�P	���,��s�~�q�����]6(G����U�D��e��o6��W�f��`�	�β���&�c���ij~Q(;�|�'>�'��7>�7b�����_F�bUgO����@�C�GB�#ϳ���;��sST�S��R7y0���)F�D+�tT�LL��eop�"|�&��zu�c����#v�=k9��=�c؃C /jvXlxVHYEB    fa00     3f0bT��ݣ�!g�00ƽ�T(��j	(���?�p�H�݃�1cD-)�1�Uh:/r�6Ҽq��%4G��n�}N�~H�rU������Qn�7)|�H�΋�*�W���3���0K���0��N�(����p��	I�?����ן����cבhTğpd�2|��KN��ܗ�N:�J�)�y�B�[�#ଂ��	q}ų������M���`�39k��`��[`9u/�(��o�����{�~�@�|�����qKb�A��9J!�^ d�/�옡�̛°z ��8!��(��� �l	�9��d00@�u���剣r�l		��?�nn$�0��	,�t 5�	ǱZ�Q���W�8=��m�CЊ�m�-%����Ɠ������C�d��	�O/�G~�g
���ɷ���P-�#�NѼ4��]��)�ˁ�1�Gv^Q�vz�Ik�8_Tز�n�̆�of�	0��|��HZK�&��R�9&��gz,�Z{���$mZ�R{b*Fg�S��
Z�����0OE�&|�UN��G��&�-��x����$s��gb��L/�@�u�]��}]\�܎�xPL*zQ�?�4"�����* 3���q�>n����C�$����CC�-�gQ*���@+%�.��@^;��S���KWd����=�1h�M�Q�����������.���A�$����B3�r��$N8�&�E\�q<�[���o�=��y��
���KЏC끤X���#����&�0gpO�Ϸ�b�R�b�$�To�p�C���+�cc(�y|��c����#���N��)�L�Z��Ӡe��4>����f�cj�rkq$"�������D�19���[����ݹH,Q�u
��,�CJ�����
�Ԛht�`�n2 �89��8�V��i�TaI�����S���KU��wS��Q�)*���C"At��K.�d�?+�z�jf7Pj���M�M��V��.�l�p1�[p�LXlxVHYEB    8096     b20��(��Y�J�h5�.��C��uu�� M���ɤ;'0Y�=u4����"����7h-4�0	�X���� ������Fe4�(�
^ek&��M���-O$g>�6�1�׆���z>�� ~�ǂ���G?}��7{���S��r�QWs��,�/gC��m#�Ǎ�.�#�{�� TY�ޗÃ�W	��q��X��*/ֹ�I��d��<V�Ӭ���T�ڿr%�.��lu��D�u�m��CG]���1��:�2���ZD��F@���P��2�d�vP\��D����~ |�!޳���qE@���\ SWj�lVȃ&����R`���M��3mh����i&�0�i��I@k-wG0w��A��B.�]\�����`�0O���9����7��9>��s���oL,��%��(F.,����o���:Og*;|�"7�ќ�s��uU`�9��E��B�Ք�ȝl�QR���5%K�ˮ�A��r{q=����Eˏd�h�ء1�|�p6V�X@��vAQ,�{�����G�i	9,��Ԍ�vZ�泩>c$~2��lA�ފ`}Ƌ)�\ŐKO��ND�U;?����U�4�ާ�ndg��4�]������
[��Nw���Jh6����e����\-!�4~L�-�Z�Z��������Ʀ^�U�yM-� �RL��f�Ft��)~6^1��om��*5�,�p)o��+L���ì�s��Dg�d59p��m�2�}VE�� �N�js��	�1��>"�2x�r�/I@�ݪ5�	l`$��v�|h�_��Ԛ|���H�]ٓ�Ñ0����S׼�p�y�=eej|��fV�O]�#�?b����������=��ɏS���d=�W��2��dmz�W��Y��/��P��zO)�ڱh�)s���5{eV"&�������M2��(�Tu�}KǉbҤ����Ը{R=��}@�{�?ttd���޵ʝ�����!H� %��(Ҙ����|'�H9G��j�@k���ID���N��<��d˟�Mk�ȮC���~�ԭ@"#/��;p����7��H��d�kJ���zռ���$��!N��닳�E��oV�q |v{a��������z��H+�w���
�wE�Γ�����0Ͱ��R#W���*��B�Z�Ȝ�8�V���%��e7��
��l8��ᩯd���9��o4-���Rߕ�z��]f�SSb��J^��q��<n��(+D
�O�q\b&nH(!�>�`x��OQ��S���>��B�:=0��.^�:�iU)f�g�&_�z72@�����S?*p�_Z��x�W���]a�.�����F��x�����ll���"�((���'$�&)�XC8�Jq������D�*���m�:2�����zG�r��#��T�
�eB%�y�_v���3�U8�Dw�S~@T������)��T���/���� �b�*C���/�5��:��c^�����cu�Ӽ�3���7�^L_a&�#zzC2�&���/LhXY<G�^� �>�W�	Z���'8�ȧ���ڄx;,Fr���z\��H��u8.-x'%�1���u/�1���<{k:g�)[8���M�  1 �w�����~)����8|�5������68�4JH4����^��M}���S�ϒ?G�3�	"3NM}���\��j��RL���tx�͏���X��b�W݋hO;<F�aLcF-~��O�K�ys1�����N�#95ד=�ǲo��b��k�quHmP;V�
nO �{��m}�DM¢y�j�A��Y����Ah�d�N�,���ܺ�+)�l9��.{�!Xր�e'BC����M��Tt�4��oc-��`6�O��Xf��#7ȳN(��o"�9���Bl������>�t�B��ύ��P|ԭ'�,
ֶ�a�������?#/����.�I �4=�̘�R%�Ɇ�A�qF�!h�u9G��"�p�����z�t������a�����Z�ce�bgv.��)�tyn"�����1ܞ
/��AN��.��Yf� �a���0��m�m!���q+$���Jc���ꪮ��j�k=Caj��3�"%r��喐�u5��ݝ��$�X|�ςٝD��SB?�|�6����q[�Mwu�B�hգ-����X� ˎ���
>r��$bb�:�?�(�U�|
���p7�D8��b�t�{v:�d��]��Q�U̹���Y^+�}�=K�1&��\J�7s'��6̄~@������gd��jԂ'$���B�S�L�?�|E�wPb�fh�����Ҽj_���b<b�-fhL4ɶ�z]������r��%�ؾ��.OP���=?0�+����Y�Am>�ro��/L�Ҋ�[H4����0ͬ���j�(���&7HJ��91��ƙhK,vNz)�g����Ӗ3b��w}b8��hU�A;���2I��r']*@���7*W�"^F+c���r��%��g���Po�y����]r��,��<!O<���0�ME��=B����@}�
=������C��Q�Q<�V����E�je�3+��<�<��0���XyQ��|�%��wMǲ�'��,����t1L��3Я�B�̆�U|�������eZ;(=AUXc�9pPƏ�߸U�)[��8�z=n�<�)"8\�h��
��B�F�&���e�b@3ҲąE�p�
JϐC�?/6m���?npmr3�3����2���:���P�lʏ/5�}��c�K�~a�5C��~N�4֞C�.mp�nB?|�ƪ�w�<���c�
�