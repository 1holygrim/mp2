XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��C��KX���4=��Ϳ��F�Z�p���k������]�ǳ�V �?�����0�u=aXЈ5��7E���x�v�`"��+��r���:�<Hy�@}��)��Y�R�:g+�2dU�#_�!I*��M��ݘlℙ�"�xhP2���C�,I ��8����1	6���Q���ƉA��:��b�E /j���C�m5��L���j�������)h�b�cw!(˜T}<�HN���C#Qy�1mVlU����H��YV�S�������z�U�ط��E��1���ߍ����bR��y���QP���Į=�b=v��8$C��Jk�+/�:�JgkP�j������L�.o�q�������r�:��������c�{��W{����������P�PXl*&g\��G���ؿ���8����J�U�~�yw�z�����e>}+�ِeT/��~���s�Qќ���"�΀����ơ�nX*
��ɷ�ތp&a�c�pNaN��"ͫ��oٌ	�o>��X�?���`�N��|#b�<����j����N.Q��L��U�>�J�z-���$Н��z�V��/O�jֳ+6���0�N�O�WȂ��cD�H'+4�P,֑�E�5*$/�����=ݘ{l5ԉ(D�1�Q~.#����B������|"k�IZ.��:���I���t<;h(�9����_�S�l9i�N�&���x)�,��P��E�1i@#�oA����L�#�Q����l �����$tŻ"+��c{h�XlxVHYEB    1a0f     9a0�����%��TR��L��|�]@����0{�V@�˳4�������#i��=�T��V�����YBbG7�prq��,�#���h�ty6�g�y�a��5�Z����4Ra����vG[��W� ኺ���'�j�W���-2�H����g�����y~M���t�9��ؚB�4H%��� oi��϶�����5�O|�p�zTx~�1�F���zйu�a�����}E�[Ϲ�4�|���#��-�n��`Y�}Ͳ��QJ:��*vfHs�A��F�C��fm0�-�J���.H*<V�^�����h�J$±�H5�����V��T	�n�!������=�{�",Ḓ{v��ro�u���F������<�l���C��).����Aj�� ��D��� '�ZI%$}�)<=�V�g#33����GnJ����)4���[� �Z'�I�����?QB����L��6T�����͋9|��vw�i���j\3Zs�F�Ԍ�h�r��p��Q���0Z�C2=&C��������d��޿ԭJ.)�r&9�3�ӣ�UnD���/"(c���r��{$�%9i��Vj�2�H�g�'�>]Q�)����K/��(~' ����uu.5[�3^շn����#R�pUC���3�Ռ�H��1��cְ&�u Uh�*������1Ȝ�0��������O�p���@�`R�y#��);¼�H��B�D�������?8��P	���2��e���i�z:bMf��'�����ΪH��]�J�"�	,S��!��4�g�F�@
�h���X�E�7'��m��2O�Z�O-�� ���.2��VN;��0X�j�d+ps� ���QH]����ZG�u�=᯿�N�4c�Ѻ;!'�@D��$�D�)T
)����6?���tl�2֙X��c˽��'��"J�f�j&�<|�B y�<��]i���z&Ǽd�2z*<�%��m����� ��6vs7�r�8��<KH��)C�oYWb+^Y�0����Ϟ�5Z_A�٘�ȵ�)�F��	I��p�>]�,�۟��xN�@�s>cC1{R&��I~+�R0ፋ���
�~��V���}d��r�N��J#�`�zn6�������G�����^	��=Ou��y�d]����PH����A��>B�C������|��W�~?���rꎿ�ʋj��Ty����b�f>��:_�[n7w�ش,����N΍`;�Y )Pe�Paj�Kt�^3�S1��޲��16`��s��{�z��E6�l@�v�n�;�[�O(KO9Λ���A�/ɩ��!��M���$'R2[Ž�jSp�uȓ��z�#Z�1�XY�u�y7�al����o~��8,;��n�sP˶v�^\���dD��Ѯ�}v��M����Z�Dyt^V|]��Q��@��9wٜ�˱'ɥ�ձ�\(����N��G����a%����ޛ�4�F��kN��c��r"�t�SaN�.��+>�=����ʶ��7�#��}��;�,�hYH�߶��q����2L�/�� $�����?,;��]䋃H+��k��p�&��߼��i���eZ]�K��4�b2�#T]����$�aV�l�	Ҧ&�Uԁ7��p8��F(��״6_�	��D�9����l_�\2}5�9��)���B��5]��Ɔ���p��@�,G ͪ�$�kH��b�!�I��ڐ��|�{H�Bh�&J��"m��m�<��-���8�
SY=��';OpǘU��E D�pf���."���b���>��h��b�Ը�G�O��(RPE:��jj��K,��#r?=�#��4��I@m�c���>��j'D�)��p��Az<%A@}w�'�_�!V$�Bq��l �
�B�f��'��rC�A�y~k��$�&�w����U��0\��Fc�E��w��+�%��g�<��*d+ڽ��i��R2�!M\N���{���6�<L�"����V /OA����Z�M�5�g�/��h��:Cv��y��]���bҖ'��e�]s�ot�W���?F����"Ae�K)Y�͎�M�!A-����X�\|�����,_bxv�5�����v��n������U3x��L�NE%X���}1�����ZM	/U��0)�ڒPO&ʇ�p�f��\s���
�fjկ�
s��e$U,��F2����;K`V�����(�AѬn�d��%:WI�)����*�	����E[���و
8k�VD�3�h���Z�6n��d��M�_�/�oܹp9�Z/y��ru^��+J��a0�{䩺)�R>��\;��T�W$��Ԑaޤ@�Fh�;���rv�����Ǌ��8��P�9��V��{m�K&�H�����#lӐ���&�:8o`��β��+WZm`��'C�a�.h"5u��=�`��!����<