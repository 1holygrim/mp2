XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��Z�W��O�өL\�"��Ќ���ۄ}ٜE��]	([0�A�]������ 	�lĳts�@���0m�ټ?)OW������T��J������xY���4���h~��:')@���z�1��$'R?����g�պ�dD���G~8h�m�M��̇��Z0�*��b�+�fx�ޖ�ǩ�vh���ˣ�{+yp�
�:�ģ���̈R!�JkK�V<���D:[�^�4��J���<��DF��a3,����� ���y����Xf�;� �^�1�B�N���1�E��m��Y�X�z�9nA >)]B����Q�֎7bhi�a�M��kۃ'1����1���i��j9l�W�َ5���Ò�h����B�Jl;y��&�h�xA_�}���o�C�u��6�Mw��9�r�#�ɶ�Z�O�wy��̙:�t`h:��8�lZ�5��dO=�ͣ�z`�j��{}P��^�(_H&f'^sT{��J�}��{�˜;.���8�]���[�ў��d-Q:ԉ�)v���/{3��d���h�n/�L<�xïy~|]�g�wK�	�}�Qf�V�f�e|��v�K��Px;�Eƫ�YBk���iȆ�csM8Q�&��X���8#fD�t��F�a#� ���`�_�49��Zh��N���ק/>C�+�bKE�j����a��~���hx�E���-�#X���&5D�4��p�~X���t�s>;��/ϒu�V�J�93A�qe���͸od�y��M�Q9��������0XlxVHYEB    fa00    2840�{�%��|@��#�ޅ@�3�ڽ�;b�5����z.�F{w0�70C���x�Ke�dj�_Ӽ��g8�Y��3YͪV8  ȀMx���'2����8Oj�6����l�C	���%]k�w���Q��yu)$gn����i���V'o� �l��^�1��T  ��	�F��[w>���V�K���4$yO؛'V��Lc�O?c.9�R��qWWlz�SY�� ���^w.���:�U���c�&�k�<��K��.V���}�ۯ'΁]����bZ�E���������+�sL�P'�@W����;���'�H6�A��Ր��)��$%�����3��b��= xI[��\�w]iP��v��ZY�v�)L<݀�����-	4�~&�*�\��&:��FȾW!7����)e��#�������b��h�e.~l������=�_�\�+.'�Zx�Bkڷ>�m�ʷRj��wj̧��=m��HAJ�c'��b���v����@�.$���1	0d���冬�����4B����Xؙ�%�<���F�	h^ v$�Y9�hVq�;��5���`�1�taf?tt��S�)�韮��I��#i�)������P8˫�>���7:q�����!��&���v֮R>���϶𨧾�R�fh�Q��Ǻ��P2�%`Om]�����)'1C�1��K�P�Οa<��l��{�1l�\*�m�`<\6�K���7M9�ۆ^��B���^��ޑ:�.ԛ�Fc��+�]��J�F/���]Ҵ�k���E����nt�0g���;�a]4�.*�v7����r�2/����("�\�t�+&�bM2~+�(a��D����������1��%|����
�����2U�N� ��/�أ������ �p^�= �ySh�&�0e��'�-U����|��/�ɠLQ���Ի�˝����υ�)2\?@(?���k�(��^J�t|��
YRC�T&kYgw���}��F�i�Y�oW�]ٮ�E���8��z��[���:ӻ���y������|P<G{��u^ee��=��1Ȅ��� �x�)j�����i�=�%h[>�W��6` j��%h�\p�r�.��n�[RL�R���[�n��r<�b��9p�:��gH�Eth���Ʌi��m��l���"��Y/�C;K�o���ϖ\����c�	���f���6���X2.!���,�t,a$k�������	�YU��������%n����`E�Bz�0�ڕ����s�����F^�g��Zv����� P�/�k�P����y�}P��u��D԰�����,��@�{�{24Y����"�rڴ���+��z�� Y�Ő~��g\�W�Y���
=�PyJ+�rKO�Zq� PF�V��9��Nx�
�~2i�����*�Q4;��'~��Gj��]����v�qQ��I��b��1r��$۾TOf8�ǻq�v�{��Z7D�u-�b��Gpp���3+�졿ۗ��k�ˉ�d/�7�GXf�d�ސq�w�`��i�X҉!���S�$9��5�}0g���
�6���Ld�Fg���Ѱς�ؑ��7���<�U(f��+Y��)X�Լ�x&��~��ŭu�Ns�ޓ�ޣM���0�t^��3��L�IȎC��ڑk�उjU�-G�ez̯
��!�RX+ͨ��@O���ć�Z�R���,��+�ޡ�쵪��x`�N2�;������V�N����k�z��3�v9��Dv�,L�Om�ƭ�"�������)K��tf^�\)�!�J	�W������j+������&�����#�@ ��0;ǡi��GK#����|faF_'�9n]hgX�v�E4}�Ӈxd�Lc�"�4���q(J�pQnjm�K�yEϽx�*�/��.��(�g����E���:����ղ��E�6�
р(?�/|o,O��Eֺ�B����i����yAȅC4�+�I%r]F^����ٴ�bR�=~,����⒣q��*'���ji ���h���M{)�_������K��9�TK�� $��H9'�T-������������dT�iE�� �Օ�<��!�p>�&�,i.r���]�9��֭��;)�@��_keR��b���GQ�Em�"�R�z|���Q���NZK(�<�a�՘؟썭Ch�ri�����f�S���F؍5�~=��5�V�d큅����ݦn�*Ѭs4]�ǅ��DK0ě��l^�*��~���5���L�B��8�_��Qxk��]O����\��4���beyv�����䤸���m��,���׍[)p�s���Fy^�S@s�0!�H��%��1X�ю�;mMx���t�f�Xd��Y�1}m������hc=��`ƫr�$��UBM�y^/9���U9��,���W��m�p�Ў5ж�j#*�h&h�^7��nc����"	�Za_{����Dt�m�}�����M��{�){��a:�sd�v�hAq����'}�X�`6)�lO炠��.�U�T�a£��'��]w��]�N=����}���3�T���IE@�6:�'�7HӞ��M˓n� � h&R�F6�DPu�]��v��Q���]�[�Y�������+t���:�7��%*�]�g :)b.	���nقz�y� k �������Cr�^h� 8��a;V`��$B�,ʨ����l7�p)~��Q]&�9,h<��+�Z��]
��ԍS�n]�I�b.�Wo�5���f�;c�v��F|J�|?f�?�5�⌫C�$֔������]1*�jU��9��h�lM>k#��A3At��hXXS����xW򪛇J�)����_�`�
��pը(�ӊ�������R�����(z#a�d�^$��*��Ms���ܮM��<Vk|�4�P�(��m���%o7��W({�S����C
�����r�Xc0�jA?G����z��2�P
�b�C �N���߬W�<�Q���Ǒڙ��9�4�����:�	o��q��Cfx)+����d���ш����9uC��i���ƍ��q2�G�^�X��:򒣰�sH��XO��qjE?����ʜ�&<?}E�p'��j�m  ��Zk���؆ށ-j�<�ܖ�������iX�o�qT[anK��W5�8���± ����������2$�T��ˢ���Q�祉:Ȓ'�a�B�D�_ J�Ky7,���Y�������|l�p8&N���u��t�<�^�4b�Q�cд�1k�[ԁ��s�������|�2��^:��P
��L���T~h]Y��W����M3�; {5�ب���A��~���h���ޤ���p�"zS8�{�X�{c�O�<]v�Β�zR��=�`�˞��D"܏�|e�m�v�$�k��K����n's�Z+z����Z�� �=
S�B����K!����g%IZ7�Ǚv2$�{{1c��v<��+D0S��%b�B�L2��M���*�&���9B�QYЙ6""U�
�#���e�nm����Q���/n��:�����<�M-�3�INZOqS%�#�M���?�D"��C v����+@��W�_T*_+X�l��?v!h�t��`�f�B�\|F���6�ߪ��6I�vf2y��]�GGq�,��m�$���|\�}ˉ�����(d��#�q�R���U��Z�u������/�6�`d *EO5�W�c�f7 &9��=m��H$�ȿ��%!�»+�ື��|P�L��b@ˊ�� �0����,s��1]���c����ɩ�08�l;�o����e3��	㾧�q#x�<;@�d	�2���`־:�֘ v���e1�p�Ra�,���M�����s����p��C��SqZ4S}H�?�XG_����yi���b!�ufp��3x�q�l4 �����Q���F���-�S��Bo���V� XQ%(�6ǣ��'J��U��5�85O.@�!iK�����)$�{���;��|����� &
�f!��k�:Гb��F�7�ھ~��.���X��u�R([�j��9;�^~�g��صƻ6y��㍾�d��(�^�SI�-�d#����J �(��/5Yb� ����4p����q�s���!��B�ϴ�s%F�~J����q���������x�D��4!��#�PA�WcM�+����\P! ^T��#!�����|C�J�� �#?�oOn�l�[�J�S,��JSi�B��|8$܎���x�B1@���.�}�j�9��pNb��أ2��%{��|����A��8?�T'N����D��E/̆ey����~U�)?1x0�Q����ب�����%_���i�4���h���V n��\������Rpf�]q��m��څg�������e�'�g�Y��C�7q��H:�3*l�p��"jֿϫ��Xm�Oǃ�)���O>@�:���5�y�6�y8�(���[�A�H�S)*wݰKe��V��K��x���<�l=������C�)	h\��7`>�Kh�#d`J߁��֛ܱp�����e>��1���_�6��)�,?����8ڥ�}CX*��_��d|�y9n��ք�{���j���4�@�S?	j4T� 8nP5�5�7�3���>4��YD�t�ʹ8���D�^ @�ھm|X�����<��@�VNQd����8������6����s� �KQ��%/�p�	n����[��9xb�E�~%�u���Zh�:QqI����{��4Թ��&ò�a_�����}����f�$u�{���$ɴ�8�f*�����.�>����m�|�<e�0����:$����c�=�]HOBQ{k��f�j0���巔���I�ȫ��XQj�+��r�ٍ]�D���������0p�]����2�LVjw��M�!��$�q���7��k�<M�4��3@0qVز���������ϡf_b��l�٦뜁I��g+q�݄ii��/��S@��ԘWx���7�F}���9soM+e���7����8+.�sa�׆��U��g����#Q�����{Y��	��8j��o�Z��uՆ����i�R.�~�8�|��ߎ�vKⵈ{G�Z�ʻ��#OT�\Pૃ# qǸb�>�4��}<.#�S�T�(�FH�;��)�Ԫ����,�9�I?غ"�w����@�!��U�V���ߔ�d�4��xF*�,8���Ѻ'��Dk��=n��xm�O޴<a���=�~�������9�c������I���Syb�ݙ�: Jf��N�ۀ�P_jG��	�kj��0o���x_�&:�%�P��|l�#Lh��|�AO���W#u�D�1}�m���]f	�����p����p-���r�_�5Z!\�y�X*h�����uˢ7b���8����G;���v�c��{��ԥs�#�[��{��0|���_���LDQ�Kc�h�K��ٰ��o5������>{Ţ��[%~�JG�G�Mp�����ouq��ۍIW:㱑���'`Z%��P=����dO������OFz����a�GTx̏2��\u�|Fz� 3Ȑ�ɓ%�-誖6F����b�Ac�#<B��Wr@�<���S(����hgBJ�BP��;�-���%�9w��&@�������i����DZ�h����kS�S�{�	���F���]�=������Ƚ����)Ȼo2��:�T���!�<���oj��K��I��+�I����j�4�la�'��	P����@����p��/z���X�(��,�t��t�M6�&�ш��XK~��޵���@/%�;I��n�4�4O�·�M$׫����t+��Z�C�'�B����\7�� �[�g��.Uss�F���:GťP��6�)��@G�5���&8G,��$|���m��x��!U�ҵ)����4y+���!�{�mݒ�^��7���\�eY�]7w��A��r1N9��Ǟ[_�\6�q�(��KolBTq5�4��*�ȉ��;����b@��X�gӨq@>����7�5ܜڕqȇk)�?��u-S���v�k�	4Y��(��G8!
��Xᐅ�}�����-�JN�a��
Z
֢�O?)Eό=─�]��
�M5t�{�b��7G,.ʷ%1�h����׺"�.�Ɋw��(�hz[�]<�짎3��/>Ѱ�bA^���!P��=�U�;�ܟ@	���@-gwy{��gS����I����ތ�=���!Μ���ȁ��Tƀ3(܆0BVjq?D��,��Ą�ڿ�Ͷ�ǜ��n��[.V���%Y1�����eYi�pbN�/UIZb�Ԇ&���h1Np_s�ꗣ�E�"'YZ���e��d���� ��%3���&`@g�AI�Wv�
��kZ�G��z?�mC��8�9Y����P%v���z�
��+=���$�����!׬mTR�M`��ILN��`�����zi���xn��%c��X��e�W�IS�KW/@8�P��\B+�T��G�cB�Q����	�V栚�E��wzZ��A�Խ��pc�,�+����L�!�H`S�H�PX%��*]_|M�C�}�u�%�򴿂�Ty�\3�+k3h.'Ւ1�h�o���in���`w_�K/YA��V�:wm�?2X4;ֹ�SE��W���h]�|�k���A֞��Ul�^���Œ��MAc�;�$�ѻ?�r����f�#�a�����9���o7)��<��BC���I��c`\��ħy��;��P~=�/�����
��&��McZ`��A���#����9)0�N�0���1֤>��D8����y�wpS�#a�d+��˂"�y^����gT�g�9+��͹�ש�D2L7�:FR����x@+W�2�9��3:����m�4Cp�վ:ktH;rݘK�Ј6�������3�������ր]F(��7�8#`T���Ԣ�IRz��]4�����zF��P��<�A�g�O�M� aL���U�!7:���@j����;Sx��+7!�R��_���1�D�V: 1Ɯ (׮�r�v�ޱXv7�|�O�����K�1?.R����HpՔ�\a� 7����ڡ�Ў�-��$�W�|5wB�02�r�ȿ>�|"�����^2��r��T�up���џ�O��pd�/��,Fl�l�q�$�ީ|8��u���Ҝ(pQAD����T}�`A!���G�����̕���C03�"����}>D�K[�lƐ��կĢN	���+�(�C��+r����J1�:�r�<�L��t[0n6M��캲��#�Vq���4mC��J��
�
�G����< �u��Q��&:ni�e���}��szv�����R��#���1��~���~��,|�yȫ�u"��$�
�mȪ"�pE��Xh����ڤ'�zA]���Wj*��aY�D�W�j��Ջ 2JjD0�'��=zU�:���L�l����"!Ø�z�X�?�9�,>��(\�(�V���b�/�j�t����ܴZ�~.&��Ff�h ��~|�*�Fg��ˋ�)�&"9E_��J����<Ĭ����{�".!�`�Ӥ=z��0^�k�J�o�{6�sU���Q�e
�y�5��L�yH[���=xq�(��V�Ra���/��x��!9��A��6QK��r?�����!��ϯJzv��&`o�8�⬣ү[�޲|�U�Mr߱d��@���soO�aI(R.:��Pat��5�_��1۶��J��p�6�Sf�U#Vr�j��YC��O�ľ/h
�x2Z'P�A����^��jJA`Bt���~]G��1g�}���}	9DfJ���(��$C�{\�Al�o���Ra������"��'�j��9������oR���dgb'�-�UA�'�x�4������x�H�yv>��Z�E�6��K2Ɏϩ/��m��&�?���،bY�$"Z<�29_�.�pw�䐡qb�,(j�*54��Ē�\%���Z�LF�];��s�2���܃M-Ln-�M~�G�������v3j�- 0F)�s�9*y;��5�� ��p��m1u"��$�,5Ƥfhb�8�	�u��CT��e���S�l��y�`ƺ!�[���`D�aY/oO���i3kzG��ϱAw�W����X)+��:�3����p�W:<�~j�#5&h���g@�u�#�0���WL������]A_�r;�wώ�C�%~m�
-gMb�<�	��/ȉ٫�1�0�*}7m*ݍ�bXY�ࣚ,�|�}�qJh�l�<)�q�]Q�y@��3����m>B_u�.I#�ҡ =����k�u7��>7�2���g^�+ÝEh`�ԭm�Rr�E �#v9���k�).QC�:+{E>�o͎\Q����:��|�K�N�i�L�+Fow%;*k�ʵI�~�:�1Ř�968�����Ԯ�0�Qς�b��y�O<S�5�;%e8P$G�Y�M]���'#%��͠��=A dC2q�:U�)|֐@���2����G��(�͝q��86�@���kG<�<2`�nW�`��#������}�V0�	,>�*����+�L����|�j˲���E�n�=)�NIoD�3���D[�H ���a0��5H|z/><�Jd�e�@e��ros9�"H�(������:�zm�}���l��<�Nǁ("uT�?�/-��~i�JM���x�J	��r��C�����ʈ}��F�ޢ��_��1Y��c���
T-˯�W�}6��w�"��|���9{�߶��Z�DZ�\��쫾�^��ގ����+".Z�Tc$�E���۷2�Λ�I��dl�&�KT+*J?��=�#y+;S,��^�H�!���-�Ҝ���l �è���{�Z��?;bU��`�&���׭Q��%��q��$��=Rj�U����_��J�H`���&�ǍBͨ���h��WE,Z�E��[\z�	��~���ȶp(>(�sM#�ӱ��?�M��2@!����@Uo�aɣ��
�W�A��bs����Q㋦�]ʓ�f٤W3G�I�x�	|3�1����j���^�Oxa�q�`��e��\��;#~���:f��t��_���Uy�Z�2nfp���|^��o+Vk�:������\�����F�¼�*`�	|�U�o���;Z��eT��n�jm#s0_G��;}O�o�&�7C;��V�2��Y���Qho�������4�v�C��)Y^�2�<sJ�+��W�,���ߴ%�Qld��mKt��?�-l��:�u��5����d[���c�Ԭ�f�����+��aεxȦ|���0�ٻ�z����a�_s����fE/�G�<�^�6U�Y�1�']b�j�t��NZ�=�#m����-L1>�Yv�Q�y�M�=@��?������n�-D �^��§z,�.�ge��w%D�!�P�q@Ӿ3?J>V��	1� �����]x�s�W����/�n�Ñ9�~�������"���u~Q�s��������5/�E�u��h��
�}[ftN�%D3�z�Gՠ��=��.����;TJ����̻!o+����+�BBVB6O-�J�1�c`�?������3�����,��}r;�e��R�Dh�k��ʞ����pX�UP� ���N��#��v)|��
dy�D���-]خbU&�Z�]����U��+:-�z�+-�M�6Ő�zG�?�W=�J�Ʃ�L��A����':�2�}�a�o�G*��GP���뚱�����
$�GF��N��3�9u��{8���4�F��4�I�:qU`1@��8�ي7~����9(��?HIw"Ӡ`\?w)�h�ZNpⴘ�$���3����a�_��Huݷ9&��.�i!��n��8P.D��;��(�95!@�iY�6�qePݡ�S7H�G���ȱ򋞒Օ����H�����tp�&�w����dO���W�r� -,����	:�z6&u��h3�~o�>L*.��ۉl��[�T�P_|(d��8g��k������^�W��h�8h�C����7��"
�"�)l��s�4�&����G�-�fXlxVHYEB    a278    15e0ꪎ�����Vs����H}�9���g5����8��[Lx�c���$���T*�ױ�o�N��r�uġ��a�>���Du$���ȥsj��l!�!��d1���6�ګ�+}{Ѵ��Ws��AK�n��������L{!��®��.]�1���4/�=	��X��hę�s���]2ujd���6I~�EC�`c��M[m�Z+�7�*�/X�o2"�o�@���qfӬ�zOZ��F�P�5Q��_�z�8�@���'�~+]�(��@�?�	�8��"�4l�d��BP��#���{�)y$et�V41n		Ϯ\)4!�_�d �6i*�&U �P��#�:��[���W�1��ŏc)M�@lZ�P	OB��5�?�<)� �П"�j��]��SAcg@�]8)�M�m򄈜B|����5DլP�����*��S9rp�r|���3I�~���~̯ h�e��e�ap��I�����v�yH���}�5f7p�z�C�y ZZ����H�,Un����.<?����2��������V�f��e�D	��G'���=-�hޯ4��h����@�>���0�)�3����/�p�-�~8Ӵ"���K����ћv@j4f-Qd
�k�&;�r��J�G���y���Gw�ϧ~�edW~`���_����~�#�IB�?�5}��7u��쨏qs�'Cc�N�>r�~Oň9�s���!�!���Z����|c�ERE#'uCl��h�آ4����ø����rZ����PtyzE�^�01#�m��5U�(�s�-dg�܃�;��K4�m�e��729:�O���D;��Kb7�����؂�^bqh����n`R��̘"C��M���G)���m(��0'����}1pF�j���M;F���/���Y����[H')J�uY�L-�g~f���|���3��5���$h���	+���\<��sw���dM�wm���5,���S��ߐ�ㄜ�0x��n9�=�����s�3Qh�L3�ŋ(��% ��b�[�x�N8q]K�ɲ����U���"\��*�F�{Ks����yo:/y��Lܷ�����H�Lm�����u�F~�w�mAF{oV�^Z�%]�p�[�P+T%G���������;�C�[�FIc�T�X$z��<����'�� ��0D��Nj78��z�	Z�g�W<���>L��u�����SAW�)�\ZEG(*�u�|�����y���)� �a\�
��{j���5�a|u_0|��=�+�^W������Tr@%k��8�v��� ��B3�B{�G=u�0��^Z�V�2QuIx�)-�R!N\�ZAa���=o�j>3� ����H�n?^�LI"5V���E$��*~�|� p�O���W		�B4���y���`�xx:�뿃�6�;_���͈STR�}����y�|�=�e�"�Vs�y`�X���'|�`[�{�Pau3���H`J5�V(1`Wp�2v�%�s�D��6�+8��Eg7�Zq+��7�WQ�!�X��j���z��3��V�B�"@�y��6���o�s.�������E��0b+67�I4�/_�A���^���h>�k$�]n�t�I�{�w�1>�-�p���#�nZ�%��ըAfj~w���%�{������x���Q<� ��|�}N�	)~��(<
0{ޫcή�Z��Q��ͤp{gW���OV;�D� E���t� �j��:���n�?�?��� �vsld��k�mt�:w�c�#%r�F�y)_�u��6�>��.�Ơ�q��}�w�@S��粸�����Y;#U܎�i�.Lb�Px~���q�<���M�G�5.�Ft,8p
;2�`�h��8;�z}���Ơ�~)듵� duH�	��_����́9G�K�1-�d]����̲ٶ�g�i�X��mWq�Q�$li�K˯�����
��E)�Yih�"���3�	�XVJ����C����N����_CM�;al�uH��n��h'�a���5IF#;�49|
��֥�9��!Yש�o����3Gq�(��)���J��*���!��3��Q}d[� ��T�'[�����_S\���|.Ӯ�M$ZE��<�Z�:6��mP��X�+�_�EZ�힩���m�a���MU��G���LvT�d�hջM�D,��9�>�ev��->X�S���.0�$���2zqp�w1��8��/��"3����$sCZ4/e�ȃER!@�n��$B��Թ�D�~,U��'���pG�b>��o����<���UkA�z6g�m,��S�28hH��(�T�*����@
r���/�5A�#� ���,3�H�K���?:�,n+y�6�u�� ��l�qH�]{:1P�x;�*xr�)6��zՓy6�\#i���4�~С]W��v���,u`�e<{,_��]�,�@S���+.Ƕ�"���:�뛃=�>�Q���5��E,�zj~!��I�d��^#�O\��Y�W.�!�a��jT�u��h1��1���?�#HW���yݓ�ò��/�&2������m@��O��>=1⬌�⇉��"�:��Sn�|��6&rv6���X?� �[Z�"�v_�|��� i�8�_��(+ í�2���{}�
������FC����?r$"t��>*��	�(#��$J
�Z��V�+]��������xu=Y Q�98jS��4Ǣ7�ib����5}�|~��x�y��'m��`RnP0���(*�C�۶fcEO����x*�QI��F%�s@P�}���.MF~� �0���h���6��j��CϦ�+��1��t���#P£b'm"��4o��*q���Vm�Ѵ8\��D{_�{�����#T�[�~ r���j2�D�	��8~8��e��}Q�E��!"j��"t���շ�`���V����(Ow�UM.��qҔ�b�M�q0G����A����1�c[O�Tm���Y�?J;���G��wO��fV�3ߕ;�j
3}D�Q��>�O��Z�"��d�{q���X�r������b5;���[(5��w/ҰS��.�tjq�,��e�k暤��WE��l���ޠ�K��ַ
�(E#�:׃2-r�ŐJ��/�j��c)m/Ga������K"! ��(qT�Y�L��@c�1�.����OEym�
�pě��(H���y:��崵�b#32¬l�Y��jC��m�^��ڹ�ћ�I� y�x��;���>��CF������0s�2}�f3�b��?^Ue���s�O�#�+��$� @0�'TKt��V��\9'��h����s�e�֎;zG3��xz3�V��l@��ϭ/�r^S�9�3��O�ڢ��_����a�]�y�SR��+�4�k���ɉ��S����*�E��q�5���m)t�m�K�QD��>�5y�t̬��h�q\����Z�}Hߕ�M����DSw����mt/��H�9�.�a4NC�d�s7��x~t�qz/�s̠���lg��d�h-����ȭx�p���F���������kՊ�#�U��L�Q+���F���C��\�
/�yҢ��
	�0*D���HI�m
XSJ+ ���6}&�-T5��r!o��tU)P!���~���V�i�H /���'3`���x�����C�r��nj'�P?��s��:�`� c0�j���q��sO>�FfOE�y���Kn��ū�[.�o�rY���to�CY�΃��:�| }��x�f�w�@\�H�{���O��`F��CLuY��\͈đ�+����F���Zz�1�������@�z��!���Koai�X��e*x0	6��j��q�J�y�������h�+�U=���f�P�"$@:r���a��nSE.���}v���l��,ÐM9,M�S�É�??e\�����*:���?���D�_7t����*q�%�[��.���'K��V��j*�+O�g$>�w��Be]����R���켖�l�9�rޕwe��ת_lH��(��,*��� ��C�y쪆zԇ?�$*g�묻�DCCSBu�3�Ri?���5�J��\��FqN�Zl��T�'ҏ��n@�+��>�)�2�o��!����Ps؍֝9�J�!<_(?Y\럥�y	,���z�	���	��q>5���3 ݷ��j�v´i^؇^�0�]��r�'���H+��r^]5�K0w/J���J5�!��b�|6fIK�k�azҡ����6.V�����-�w��#S��L�:%�ø��bN<>v�Yۚ���������,S����m��O Bpĵ��x�-_8΅��aػ2[�|��!u4�����N����Y�����,�q�vckP�V��䂥�Jji�7�����1B�^�����P)Е\|:����6f���F �I�]�aZ��"������P��E�C)S��\&L�g����N�5��5�,6��V���mD�N�f������tQp��/I�E)����}��/��z~Chn�Y��Ϩ����v.p��y���d�n��͛
��V�N)��sR��-�����A
pȒ��L��Kr6��d���Y�(v�:��L�Hq�ƿEt���,����Gu��E�vĚ�	3�Ϸ�at��=��-�ծe�*��RD���j3E�j~uh��jOV<���7���!��Px��4�����	�ޡZ����t~q�v�=�Z�P�fK�օ�sX��Y�a��J�&t��k�F�#�4'˛CD���0#N��e6�Q^$>)�j�*0���֠㮙���V}>@��u��2�KQ�)Y Bf4�bЎ_.d"�.j�$��9R��{��xͫ(E��퀳Bu��o)=lj$Dk��
Uܫ�\��Ѱ�8�3uQ��v�㥪y�/U������]QF�=½;ՂG004���Զc4�l�zO��O���ŗ��rY��n��E�G�"+0#����2�����&i��e[�~;�6������6}�,F�8̦P ��9��B�
��9���5� �0���_J���6\���+���I�&ا�,�g��Jow|���1����5���VH�~�9a꫖�	w�;�C���xHp
�m��tRTVկ�]�`W.��?0wRt��̅]M"M�M��XD���n�v�~�Ԡ#������D�&O(�nh[M�a�O૦l�6XY����v��j�zR��~��$�z�sy
/�YY$�o���o�u.����p1R�/�r!�4����U��L$�	�/��*��gފ�0�7Fq��������Qw ��(U$�K]*�QT�5�P��o҇�d�@��a:]��q�<Ԇ���V���þw���g_q`���yi�'Z�:�onm�r*��:�+�O�ߦ+Zi�P� ]�}tȔ���?W�a@����\tf�ya7X`�)=R��j��qp6-�(�<�)�1�;����!kNa��4��p��$t[JD&6��(�j'��!�5	�f�͹���6G3�N]LO��/iw�D�T^ᎌ�jkC���V�9��D�n�o��_�