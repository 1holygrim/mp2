XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���<j��0�)E.�ic����:���F�*o˱��p���}Y�f澞�j���"��5�����ZuW�K�a��­��0t��zz�3�6Gɶ��i��z�c��!���s�������攑�Z���!?�Um߸Sv&� =�^��k��@�ԡ0������팺1H]���=^8;�	 ��K{�Zd�0����� n���k�����:�n�#���[�'��h-�[ �r��
�L����N��������l/M�+ݣz;]���l�����G�n^m�Z�Yj���z����:0b\���y�r�Տ�yF��/����~�E�#$3�b�[�T����k�s��82"�Ѡ����B3U~����r)m�&]��R�Hu @fQ=�^�Ӄ��;�#�ؠ'J ��1QQ�0�|�ӸK�:�1z\�r���w�б�t����f�QJa�(Ps�xO�i��g6���;k�
++Ñ^]�ln�8�,kq - "u�:��9I�P�^FW�n�l��P-�UW�ۈ��Տ�Sۆ�F>�φj����~'!��L<�\�<��w��K'�⓻�'r���[JG|SK��lB$��}Dx�u�����h��B����h�ڔ_`N��'�ɺ2śɅԵ�`ˑ\5��غn��΢n���=6��0��Q���Ӱ���^����UeB�5)-���`�W���d��@���'���0qq�r��r�ީ��.��I:P�#�ݚw� ��կ6,5�9&�B�P�D*�)>�34��In��nXlxVHYEB    3e93    10b0R�Ev�`_o!�ע�΃�x'L�L����2��rq`Ȯm��'�vPLM딍υ�ܑ ��F����"yBU������K���n�;�%�fZ��nR�B�ͬB����\�dBpL�9�.�`����mG���<�d�iLb$���D�)���>�Y�WW"=�]DD�jJ��Pϋ�)��d���*˚���<&�vCⷛ�.�I2`Hme���}�jE�qb��ծz�q##�_>6�h�%����#��>�"v�*x�!-�p�ؗ�C��8�,3�F]u�W��aV����tƩ\[2�.x�n�����b!�!��b�f��
���HԊ�����!6IֻG�]����7@�c�o�T�=[1�����H�n���,���T�^�����+��sX"�Ԏ�<���G����za��~�)�� �Dx���кD&��O��3�}��S������/Uz,�X����ȳ�[��C��&�7�����V��L2��x������J������kI�`e`nPP)B�������������oJ�љZ�f	6I/�5u�O	T7�
y\�Q�U���1X��mzm/�m%U)����N2�63w�������k�9&�U}�e*'?9��00J���1}��x��JƂUe����,w<W��F}�;�=�f���1^ZyLk�;��p2F.:��F�3��e��X%fwu�x�����E�L��&l�I�m�Z�"��B�egl���!>N7CUKH�F��j?ˤ4J-��nl��Fct=�o�e��9)<ol@c����g�2���[ItJ�F���NH~�bt�$�4u��J��<(�A���{m_�j;�tɊ5ay)
���}�Wf�TwG2�s��˥I��ߐ&�0Bw�u�l �:K�ͥH(h��(�#şZ$�r��k�l������[��0-<[���;��3��SFHκ�F�3��S�2�0���뷟�L;�VEhL��>m��ɟ�u,�R�HB�$�a�����abhɨ(N ��Pv�5T�+��b��X�0Gh�=�����O�H���\�I�s؇s�)G�))��, ݬ�Ȋ~%?�㞾|/��r�'f�g�"�ġH�*��|a�/�(���bh�h��°f����D<D�`��N	��(��OĿ�\�f�V?�ڹd@�k�A//,�1� G3w��ֈ�e�һk�PS�/�Z��^�'��Qp��J��9`���V���i�� ��#Y{�����o:��g���qγ�R-	1+j�u���Y�<b�" ���2_Ij��Tba�����}�X%d�u�5�2��,�K��쬏�����3�c�ʹ�������%��&��7�N�
���9l;��qkA��{�5��&�h�0KN�p�a	�!ur��\ka�m)������8C��%\�d ��@;G&l\�a`*�y�Z�n�n�F ��17��N8A��i�8�p��<x�̿7��0� l�|?02�����C��_��.9^t�C�MWI!EP��;�J�3[e��BAYZ���5$a������k�/�h����<B?2�f�G����ƅU�3䅩3w��=��f9{0//}�F��� ��lu
�ra����IY��Oߘ�(]`��l�0���M�?��y6���N�I�	='>�&ӧV F	<�	:��;e�����H�{�C;�f����y԰�j���lu�������o����:!KG0�����i�G�1�ȓH+����pHVxܧk٪���v��wvB�Jg��Wcj�$N'
�6����1��hψ
�r.�	6y�}<��]�m��/���e��u"s�n�P��v�K�y8�ًp�b��/O��/KO���� j\.��h�%���Ȅ�P<K�>�-�� I�]N�M�Gf�i�%��.�z0m��L��\�z�ְ�.J ���_�R�? TiM8!�Be4��+��k�ǩ����$~Ig�D�E�:�4��K����
ҙe:�93ֽ�=�d�����2y����9�a�#�m�����<����a�RO�jIJ}� �M+�'��I�Z)Բh�WSXO#��0��P��e��w����0�%1�w���@�]S�z�[�*��MP����m���ՠ���Ң߼��-��!��������[�J"T�F���߉�̵YrIG��,`����>'a&��/�d�~;}�ռ�m�L���T�� ���@,��=����i�遽d�R򎪿�!�U3��u� ��N�u�B�ċ���+�1�x
OI��N� c�W�Wq����^� n����P�����y�\0�-n�����h5�8�u#��&�am����@C��j��ԃ7�\8��.�O��+�:pO��mːD9D�!�@������s+c��X��t����2�*!j��beAW����4D�ಧ!��L}W�r6��W�F�6V��"�Ap������ɝ���������v�]XK�D��}����;]�c���ǥ��i�X�B+�S��
b\��~�(��8�,�ĦZ�|;��
'��ŀ<����U9]*��'��Ȁs�+�-��7ǔ������X����X�&��)4T����n.�!�џm�^����'��zDBCYz�۟�1��:���=n�n��!�:���z�L��1w�Ƣ8&��'�#�$8��"�e+�R�Ҭ[�^����-�Ñˁ�
�Z侟șٹ�����Xè�w�y��G�2�W\CQn` �A�u7��:o����I̵�Ν������'�L�a2�}�^��S������ �{����Ipe<�CB�̙��Qe{�2���(���i��3�y�b��j*���d��G�fG�	��0�.m��n�glv�hyE�,�ũ��]�Y��g�n�XUmt;��/��m�ϐ~s�}B/g��}d��V��H�
���t�+ d������t�"�Xo�z)�sջ�p���_��V6�0%���A�3	�Ľ�0�`�p�$q��q�4�ߡ��C-d{��=�>;�s}�]��]�����>�/�X�"�� ��^Z_��.�����ʇ0��w������p�n�Vů3)��1�[_ v��g���F�y�q�>�]�|�bѝ4À�&(�t��T���
��&�|e�uj�@��֌ܔ̔&��dǤ|���{�y+�N�:f\�c��X��53D՝`�~�O^l�� ���X>L��J�z��%#C�m��x\f ��M�t�|Z��&����<��W�)������t�:&���Tynm{�����@�EGN��na�}��;�;S�e*�q�(<%�z<1��X��q�D�:�nY�����߳�kkLf����>}�q��rЫ�vx�5��>�	�tw�9l���P�澴����7�y�`�o��C��Œ]	�^������D�}�����s��U����`�t`�|�=~S�,-��<\��G���yE���DB
+n�8W������ڜ���I�����=�Yڑ�%fKDdOx�Zc(�)v!�h�[-�u���v�c[[�R�5��x���W�&��	�X�����5��Ӷ�Kl��X܍B!��<OZ�h��>��DcqP��Ǔqt,���X�5�P��|ں�4�e�P�د�a	8�eX�ay>��� ���Fy��z���p/�yMm��#Fc#Tr�©$�+��Oo@c��ڥV�b�r"�u����,��n����I�:���j��k���4j�cj!oV��l�)�x�w�0���X���P� �AW`d������c��[�r���_�}}>�Zr�c�=�8����d�^�ttC�1�w|%<~�m��&�r�f�l��|(��y�}E/ؼDc|����}�<B���)y�p�Ӱ�6�Y�$������a�g�
2�"&c�N�����h"���kW���̮�"K���G�%����������^�dN�����F�S�1!0Π�ގZ:��"�ݖ	�9p>-e� yH�t��p��搈nЋEgQ��Q�5Չ&d�dֵ��ۀ�[�֓�#��[��>��44|kK"�f�� �bEI��v�A�b� �D�ޜV8��Q���	�1�A��ٮ���ye�R�0�0�� ����vV(�C�e�ؑ��_���7�Sʒd�yD����ѽ��XH�� ĵ���GXzw��ka���Ir�wP�R>!�