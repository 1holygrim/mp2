XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���T�2�A�	I��jQ�=������`���L��"�{�-����%�ǐ�;%�B�-�l^�	:jb�d5N���O�E��C���C��ap;���'46�g���y������_�l��3P��	4e�D�*ѷFLd�Zt�v���_��=��e\�݊d;A����ޑ�ud��n�4�^��iڠ�TB5�IJ:vž�:�
����#��n���.����U� �OU�nv)oP	%�  C�;E���*{��J���u�����(�l���u��FJ7 �-�0�IJ�E��sבW�z��R�6qGn�L�2?ͤ8���\�Zc`D[po�ɮy�q�~Ē<mr����NO
�����v�D᧰�������3m$h���f]�;���/��	����<'b_�@�S��e>���S�mꡍ�����d���S�R��)tUC>>��s�,!xH��q��N?�����J@�ǌ���w(��[��M��Ƨ����]~�0����l��n����9e�=~��Ύ�LFqQNxZ�/
8Iݼ�u>F��V�)9u�� ��ݪ��A��I�T,�5c�K��'��%?3�A:�9���+�+�K=E���F�n���N� �%uy3�.�R_T�s�Tiy��P �����Z�	�˄@���/E�؄(���\�'s]
��@��"�5�)ڄ�Kٙ���mRl	�۴�Y�&�`DGyA�T�����EL�<3�g�zl�����4Y���|�|�􅩽޵���;�XlxVHYEB    6315    1790�7�"_���4�L����g������#�e�ƴo�b��'sy/�/Wp(WbUE�QY`��	f���=���߼�����3��C�x7���Og�����2��X�֮�W��W��`.�r�W�U�)�<���W�s��1	�F�T�4JF��nfY0���٠�V	�'��xpzw�����q�e��')��*l~ȁ��(��ʕ���B*���"UL��)���h
�~5����1K����M�=�J�zA'a����C1��J�o�_�l؟�3�d_��$.T���Q_�ON��o�wT�K��d�/�1�}a�	�s�P�7���:ӨE�A��8�eV�k�W�<��詌�iZ6>xs�_�7�%e�g���`����Z�⠑4��A����g�|��!"�p��G�X��l������m�D*��&l���OQ��p�z���R��� Y�!eq?��)T)�?������wg�Y��Q���G��Ի��4_V�=K�j���K��� 	���ȓ8&A}����	�� �Dд����b�mr�i'�,�|k=U']��u���x��Yrb��pT�@r����jbj*����,�����w��@#�iL���,q釫=�wD�*��������Fc�ŷ�L���Ch�����Tt�`���W�&@i��H�#�Ŕͱ}� �!}p�����e^�R=�R#�� i���	&s�xh�t�>�|���>*�Dn� �����!���P�łc���ID����\v�y25Y��Fi������]'��=Ij�ZdK-$���z���
�����X�Ƶ��VC`�`���7l	\U��W8&$`�����>�,�a��֮�Ýs���:"S?v�����&�(�8]��#Tv�v������&U*@]���_V�'��.
¸M�Dud9�?s!��\Y�g�fǌ6��o]O��0���\P������$�)�3
�8Ŷ��[y��7������^"��*�\���h�P=96�!-iE�?=z�J {�g���lz�1Vv�����f=��I��w�~�Y��˱�_��K	U���rrX���̞�	�8��9f�E�������]��l�1K%���W��`�i�7!�T�SV
vo�T-��Ĩ`����2�a�DmE<��SŻ��c���E��9����Lװ�퀮���H� `��\x�ed��-mt���h��U�~)��\;[�n�� ��[J���Z���<G�sVPtP�z�~���&�����H&ll�U׆�K�(_�����_g �OP+Бy?�+�g�5��T0�+�+��XNj�z��LΛC����.��7����Xv3�WN閂+��\ٴ&�j	�|���Pj�3a���}4#:�d�P���v����0����&-PЇ�B�}��<�� 5�X�x@ߕw�t���6��6�,���CF���������42��������Vb�}/<P{��󄬎"�F�$$��y��	�L��(��x���� k���'��SڡأZ]|��X΍y� ���Q�Ju{��)U�P��:T�뗪�b\�� �U�P����i�eD��Iz|N�4���(���F���;z'b��6���؊��&� �D��MoEct�|D�	�+�H�e1c�Bj�s�k����#�	�����%׶�g���P�f_�G}eb��d��,��xMO._6q+2�W����y�����_�;l��%s��2�B�Q㪮D�'�_�zY��)7Ћ3��Zzq�.�=�!M�EUEa2�L.&��(��!��rӨ.Ϧ�Ӎ\��e����-U�-�Rd��������/D+��S�{��A�e��u:UH���u�bL�:@�$�ֽ�bܟi��v��{ݕ�ۀi��Q�frT@w����-�N:�r5	b�B�g������[A-j�'
����M݇wn"1�]("��5��\h��b��^hwAi]��V����}�d^>��CQ�&�4�옷�$VD@�2f��~��yZ�B!��Ӎo):�#/w����		��=��ӈ���ԋ�{.�m���_{���z-�3�0�MuaN`�JN�mT�w7Ss��Qš2���"�M���e;���V�y�-AM㙍��0� ��&���H ����F:#���'��xV��Q��
��>�R�bp�\=�����rҺt���R���^�+4�t�¾cfrC<�W"e�~�I=����L*[���A],֍3��5�U��r��$:�!�X�\E\J'�]�c���>�
p����kSV�Y���I3q�?���39Ҁ�D�����f�U�����k.�0����X�)��Ϡ�N-=u�����&�i2vE�b��1� 3�C����lEb�L;�,�R����K�k/'�(�_��z[M��M��-�����2w�YE4޴���V����mB|��[_�`���Ow��/�̑�Y9��ӕ!+kjft)��Y���}K�
���jD��|
|�F��3c�������le>3-��է����mS�<�PR��V|H��,A�;�����6�Np�qON��_'����w�*�*��?Ao$XF��Q�(z�ʿTpې�
@���Z�_L��.h8�Ql���.�h^}�/�J!R��flz��J�w�ԃT����- N��)MoLW�V�w�R׀r͡FFs���cOr�v��oº�M`�^�j��s�w���<a��l$�;�>��H@Q{�.E�|�-�o*p���3�;�����\�]���|2�2�Wx @
��ؙ�V(�9-�oSbۘ����� �;b�ltjM�o&��{{���Q�^�#�v�Yߌ��+i}`3�-�Sp�̊ ���5#v(��eR�۸��})Ò���+!�C�vfTrG�w+M�k�?Lt��o3(bNf�*,�:^U4�z}�:M�,��w�:9�"u��Dirm�0��2�n!�놸y�3zM[ 4�dx�A��C���Q�8m�SM@���{>�Kq�t�ՃB�E��S�����]����f�����HTi�ٵtu���t⁪>�Gi�B����4�j��vx���&�E��1�$ *Y�F�n?L����pAc�!�/�?���#�4O
��țQ�E��x��QƍP��R�w$�<���?������+�>,�Edg��,cX֝p!�o�P�	�@�1���M>K�I�;]I��q��z��0f�'�a�<6���C�3%a�Pi7��Snzy� 5���}��4�«r3}P�����n�[��{N����7�NDB C|K��w���jS�]�l99}�r��]@;�=�MT׽�tU��9Ƙx	��D�३��"���R��u���ߏo�	u��'P]����i����=�L]G�t��ׯ�(-�<� �ms��T�)����p��Q�ǜ?����M(b���	J��}��~���ѝ��F��/�=��P�%���b�R��^%m�P�e�ϻ���5�s��@�]�}JsЗ�0�b��]ہ�93|�)�Y�+��>�/O��|�{w{vs�QL�rp�*B>�e���[y�E<�tr���.GB����I�U��b��ö�/kݕ1qp�qO��"�" )�xI*���Ԝ��[���F,�+�X
�u��!q-���vk}�Xb�y�x���Kuԥ�[��o�>��6��z>�xT�G�g�eP�����Q��yH�7�x|����ռf,��Y��w�fP@�٧[�,�"ݟg��tm�+G�͝;9}S�,dP!2�j�[��k���y��zq	����JH��D��D�$m�8���F�@`�?�J�ˬ�H���$�O8t�y>^���
�وΞin��z_�ic��N�us��-9�MI)��XZ���i[��$��-+X�UeEq0�������N�%}!��<=�GZ�0�2v{��4�����o�?
Ɨhv�@"Т,U�,�ZK�/��"��Mx�t��ց��կ9�FC�He?��q�l��D_�,FP��8_ʆSxݹHAs�Ov�����a��v\��i�D�>z�߰��8m�y�A�ۨ��r*�=�?ye��4�����'մ�-ƶ� ]�,A�F� �<Ѕ��L�R|ÑP������ȸ�K�.9u'�����*m�7�ZKqNy�7�&T���r�7n�zw��*NN,�v
��s�w��{%�ߥ��Iټ�XV�C�T�V+�F� �669lq_]�y����!J0�CB��D���s���h2��Z�I����[n��]�����`��7��V�w��l��eG��/�a�	�O�q�����ո=�&k�p�v�ӡ_C_�@�����?���F�2��p���Q�P5�4h>��ê�~���D[Đ��M���~����N.�kձW�<�~bG�#_����2`�$���9�\
��)E\��z�U��,J\�,p�3/�QQ��\��hR�l�p�%Z�J��8�pa�9ub�J���^����?�q�I��>��Հ�ʵ��fñȬ;YB栍�|d�vN�oa���ї ��m>)������&d�������+�LҊ@fz�"�D3(��t+@�eܦ�9o��'`�DQN:��L8+�i��S��.�oC&U{�-d�<��Z�H/Ǣ�\a�(\gn��Z�:*��ð�oXK�ī��E�'�h�D@��['NX���z����5�}��-��e�1��GBg�P��~7E��,ý'���7[�� R~7^O�|������8	uD����;u�7p��U��v�s�Q$�k)�7�$AOe��/�w"!	]}Q|Ћ�6�����A�&�TR?�!Ly7��I�Q�����,��WTO�Qx��T��pW[-10�5���\Ι���$�ޚ�V���-���!UL"㜿��r>�݃a#�c��EJ`W�s_�[��%��Cv�MP�}E�	~�!�1�U̂]m��VG�o|=ɳl�&��Z�'$�)`�r���WN=������)��1ҁ��zn{�
�?6H�P|(
�)t� *���""3]��_��ܿq��-�Ǣ��U�e����[=��}��W�fm�D�-�6O��}���9}�%X������;=:��R�m�&��>�Ҫ��?p�I��c .pJQ��@�#���^���'���� OɄm�����썙�=���-�`[ 4��&�5�jHy�T�p:�%֑v��>�M��mv��+S�9�}�'�^�vKsdfO(-EALصSl���f�	n����C���XtY��.�q�{�˙�}�j��h$خ��L�r�"H\��+�ͮѷ|9z��ź%�pg�[�-���G��v��]w�� R���4��.OkQJ�2�s�u���8�sD��+�BỨOK���'nlB�ypl�v���|�bu$�6��:�-��UE|A��p|�:���bR��MB�6��h�/��'����0�K� �x�]�C00��a����?����Z$e�Z�xw5hN��"��g����2F��~)�_�6��N�J7�vՏ����b�e�[}�ms�בZM'�Ƙ��.jֲ�5��x~y�%���w���`(͚7S<1�K�����͍�aRegI;��ˠ#��_���/�3��7@���A����� ��^�l��:�'\�A�J�A��;���z�� ���H�x1l��Y�2��DƗ0���l�݆ŵ��e�{��`^	��>���޹A��Ca�q\�h���S��Yw\��2��D��I��d�V.��FCF�j3�d��?j��5�_R+�W�ӌ��݆l�7����W�,v�0�tC����1kl�gvr:��YjL2���.�H�l�%�W#>-���٥Y�q�z*��)H��(/w��C+?�#B�}2A�@p��tay�pO�a�U#����:y��9O�@�e�����M��~m��-�r�