XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd������G3[�Vh����#뛣D�d���w(Cq ȼ�9^!?x� ۢr�c� ֭PR�r�>Y`�����b.rV������S��� l�װ-!��N����w�m��l�#J9r}V���$��WI�]3) ��V����m�k��kLtxT",�R�I{��Ex4�)����uD"����Ō�(蟴����ak�_���o�z�Řb4���<�H�($<
XNr�'t���ۘ1=�ӆY�kE�����Q�c���V�5�Z�bSzq��[U>&�G���c#��S�;�Z�A��1������	��Fs��I��δ��c&�/l'	�~��V�S�o�~�7?��0�` ���
��=�*$K���_$|���C���Nt�8 �%���&��id#t<�P����u ��ds�{E�(�l�]�QS!�〠X%����N&t�>�Ix淯u�!T�|{8��T�΃�Z�T���'ڃs�Ǹ�Q{��U�:7�7�ɯ�=�3��mx���L�e;h辙�~������re}'��h���)�y��A�,<1�[<�u���@H݂��!�mXݭ��74!����%�������x)�m�������U��;juvX���\�	���WR��E>^�`�EDQ�5`����c��(*���!\�w��?:[=�Or�W#�-�1��Zd*�〬n�XJ=�����Zq��B�h�	���72�7p�HJ�������P�tIk�g-�:���'�
1���etc�XlxVHYEB    39de    1170.�} p
�$oȕ���P�k��t4��[�6�*m�(=Zw��&�?�./�%��<�q��^�}*��"O3d��9���^���6�|[�|�@L���'����m��������)�V]�75w�ߑ�Ι�oO$������A�����SQ�Ȗ�Zw0��r�5f�FM��?�	7�km�k��5w�����t1 *Pu-�h":�v�u���D���UI���J
��	q�N���6��5��,3��K��RPǢ�W.	�|�
%3?2m��GF�j�}Uo�b�eX� (�l5g%D��>��5Kuh�z|4UVxn�VB�e���/��8�EHv��S�
��iس񦽱 aҡ��
��V�!���Sk"ȇ����I��[.�9O4*��w�_O>~١��	��4�Ć�B�c"�,YB;�E�,V���R�u,���� O�'U���C��B�5�6�bm0� (ˍ��bL���f<:�S�Zôy��޹5ٛ���У^l$�n�"'�6zŃ�Y|(�L����A�گ7W����5����z	���hO�X_>�O�Y�Z��9���v�s�=o[�BV�0�wG9�f�8�y>D��҂z�Խx��#��z%�gq��%��՘��t���'��&}p�@�����c�����>��9S�;�ӐW�=k��HuY�'ˠ2�b�TR�f���M�u(\H���^�9.�1���a�?p��G�C���8;a��XB�_}d2�>#�q�c,��ӆq�U�t��<���YՆH��j_����y����=3��!E}jp�m�&�,_�cOֿ-�a� ;V��t!�i���6���ܜ"\a2�"�I�������T���@M�;�a�,p�J���j���G��=>��a�өò�M�o�ٽ삺�^1Zj����3.��s#��ˇֈ��i��/�r��b��݇����^�	����L^�#��B�F�9B_b{����|�'m{������@8W���D#}HdӼ̨2bc���#-���ͳ��?��q~H����y�"�t�	&��J
����5�b �7����N'�B� 	��&C�
z��O��͑_�y:�8��ߤ7	�>lt��q�Z�cUF�K�p�\)�0؟M�(��7�P�8��j5���n2�b��635+c(� �ǎ���ww��:,Q���c_m��'Sh���Sb(��2By��A����p�B}db�K~/ׄ
�d_U�1a�˶��_�}��i����Ѥ�M�'W�	����������9�c�b�</�"��!���P�Ppw"�"��Q;�U!�C+²ٸcPw�?Z:���G��C����~K��ή���%�?�ITW�$����y����8��DPV3 �W��8 Ư����9�O�#̣�.�x��=��ƫ0w��[ڻ�NP��l���D4����r}x����OO_It	#�Ɓ)t�t����eO"YK{s@'B�/5�ť���;	�R���WYX�[�es�Y�ݔh�R=��-I3l��C�##CY4�=�z�ɱ[��'|��v+����B3N��k���	E߶Q�+� �d���U��Za��.;rcƚ`�B�R���bD�I^i~��S3p�<64�S��LtK��&� �#f�h�94�@-���gxV)T��'�Nuv@v�^�*�7�|�0D��T�����#��t���DȨ�/s6�-(%ҙ�����E��=��7�*�P���>p�n����f��{zA�0e��>)G8�XAZ5U��)�<�!��o~�Kj�k�wԞ4�dL��U"�{G�������u �@l��rA-u�(�WԘ��ĥ��B�z�{�nMt%���Gh,$��*MuG�k�3�-GL7n4Hѯf8�U�Xb����c	�G�;P��t�+�ǁq����FYChfꁤr�6.^�"A���-�e:u�x"h�F���`��м܄5���d��&�+�[�{�HX�S$���<��z�_�땓�V��W(4�7�#�Y��{�L�qeDڒf���|<�Siơu׃?���--ABM�j�k��=ɶV��$X��H���o��S�Jm� {��������x��,�(_��WBr˸�*�v�S��˹�dZ1_6���4w��,�%�q5���)⚿rN���3+�rH������J��w͑��xDt����X��P/�Rdxi+�O�5?���*ԁh�H��|0��{��g+@6��ӵ�]�<�~?Ȯf'�Es�#�(eV���K$�j�\)ս5,Sh6t��U,�ȗ�Ua�U�E�H��U���G×��O�s]�+�|ԉ{	�I�+7�2�E���~��ܻzaD�"���HV��#�~��:M�
��6#�Y�B��!�6�{�������d�2�N��J��$��P����Q�h�r�q[�C�|][E����䅋��W�����st_=�<����	�*q���OO0����c�K.�4���X��5�hO�[��Xy�>�~g�\Ů��w����L@-�� �ӧ��5Љ���j�c���e2�튞l;0D�M����=�?��V_���.����I2����(�<�/���դ��C��Cx�u����6��X�L�x(cҕ��x�\z<�M4@���ѻ�Jt����$�Gz�,o��o�0R�5M�j�`��jV�&aነ�,%��F��ᡍW���iR��4$#��3��8�?;y�_)���<�`>�j)"���_�`�b���� �g/)L���������.hɋ�@X���e�A4x#�H��1]����RK�	�ޥIm/%��E�]�NK�P��h�(�؞p�aNx� ŕ@�d�:x�E����~%-ɋl"+.�YB��d�VW�\kn�xQi��uq���R� ��šh�j!~�)*2T���6��,��ЋѼ�J��jh���j� �UD>���\t�ĥ�����4�<��]��7�KL�,�a�O�"�@�؇`w�RԊ��$l���LҦ��(����'�k8��h��r��*���߆��p�Q[��r����1�բ���n��A�N �z{�"�؀�GO�G��O����C���{�>K�.|Q�-�@�/��n*��:k?����(
�,�j��,.jrK`�|���� ���L3�)0C�m	`�a���wF\}H�����Rm�B�;G�w#���e�HI���X`81���S恚?�C��z ������ReE\�og(l��39��!���b7g�O�����9���Uh�z��h��8���C��H�-�*�W����B��lt8T�+���R�@	��T����]v˾��OD��=X����g�� ��F��`Z�������8��p���G�룾�1�Л�G�K,&W�߿��!����4�9�+mp�u{�#�SF�i�Ք���й���ޏ�T[	�z�i��*w`�F��$�B�{40�a6�}��݄L���)�vGtz�i����URAK���cg���R��A�XG��󔄾$ʙ���V��M<�t��<�q����[�O��L[7�����"e�0��1h>����0�؉$
L�w`Ɖ!�N��H�Z8�Έ��:?@X����r̯q}�9�ԅ�N&��e��B����ʾ��N=��6U����mF�i����]�ĝZ����c��O�b��ߍr����a�i�췞��W��ݡPFM�x��
�`P�=�0I�}��u�x�2��37�����`�<���xd�j���M�x�=.Tt$Æ�rpga���dT��.S
J���jJl�ٮ��P[c����gA�iqd��orMF�����GI�p����k�����d��U�+����dU�(���㲀�6�%��w���5��E\���ʸ�aE��ֺn�+t���O�
�4�̶����q�� �w�A2ɇ�������PI43�%!#h��g�te�¾N��ZT�h}����b�5�b��h�[ϟf񁘐ݏ�i�yT��0�X׶���};���Q��'�*Wo}�_X��5�����
)!���J�x'��s�Q& �rȌ%?�x�H�s����m��#�iY"�zK�$~n��G"D��B�<�w6�UV�%��r\�a4�(C��F~$7W�AmlrS��s4��ܛ��zs'7��HӚ݁��"��$E����^��7�`H��m6^	�v����Io���4JB����=_�Cm�X姛�W �n�- �>�#�|�9�����U`4'C�+�8Z+���ޣU�.��9$�Hzl��6}�,D49�8=@���<�uAӌ�5�\��Ɯ�\O�Gĉ˷^���FF6�-j�*��@K��0/T���oFH��H��L#���<~ۮ.R-=)�ժ��ap�v�z:�"խ�إ�