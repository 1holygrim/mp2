XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����@�CYn@Ǎć%��h�n��A�b�d����ܗ>VEso�c
���W��������
rkٺj����3"�[�^��5@�cS~�+YHF/�تk|��l\Q��-Z���f���:'�����������d��

�	��^Z��#�C����UwAL��%ԞzS]*$!źkw��^�����Z|�CZ2���o�ޅ3eݽ05�J����iB�tE���&W��[�A�2�>G�к[��뭁�_�Pz��#$>�Y�����O��fI��{�G/��6�^�nl��[�Kv������Єr	�n����A��|FK�t �"zY�eǍ1�q�0Ė:��u;|9��� ����[q���w=YFefݲ-��3?�^�]�W�UP���D��J�Zgq�1�
!�����e�0����;
5Ɯ|�p%n��⏁����$�����W�-�q*tǶ��Ms���s�	 ������0z��~�V\��������2T#��L\��{��rf�3�+��x[�	�W�O�價�!A�ŏ�*��������af�O��`;���U�.�$���@�);g� ��Ͱo� vzO� �KI*82�ǽ�Q�Ky�Q�O�wl2���9Q
�-z+c]�`ٟ�⸅�r�64��]���WH�L�[�OG����i�o��z:����7g�A=��Y��@�<_���G�����v_I���l���K)�>����FP�("v��lfoc_�<���hW��7���m�K�XlxVHYEB    2a14     b002%����ʢ|�h� Q�����c��J��QIW&�>�#�y(�;{�M!Y{v�QU9戩5�e���aS�G���7u4�-{�nq�م٘O�B!�� ����u��G�@U��9��@۲�J"�`���n䌻q�%95�JD��l����[��Z�1�u�C՘Ձi�]p�`��o��44^>�����;1@�bV��ߖ��쏀ڵf+�
ʊb��!3�a�CY��kC�-�Ȧ�������+];e� ����?+8n(�z%�0���8ɷ�p~�����E�w0%(A����\	f�GI뢱I�yc����C�����r�?�Y����rΜ0��ʌv�}q2Ԩg�Zl�:\L�ٰ�m�}eK��&"�4�&����9�[A�3�C43|82���h��sJ�5R����>a*�R�z'fk
J��2�o�
��E���ܫ9I�~O���1��)��As%��=�W��t�&M�6={}:[�)H�3&�R<kC@	�%8������;��i�`�k�x�{�B��ʹ�̵v6��#��žПx��Qn��|��Vjc�z_�	����/f�8� 	�#����8RR��@X�w�y��(�ky���
1���b�` $��6�s��g�TJӼ�6�iR3Wi��$=�o]�U&�6̸(6��vTۙ��:��
�:��&��z�.7�]���� �}�'k���ўvd@E:h�1:��7jk9�o����g����腕V=�`��`�ry_F-£�9Ptm�ի�7﵎�+�LV"(�NU������*zҐ���f+��H(	Mާ-�A1D$��I/�U�+b��
��O� ^�^�� �0�}I$7
�_g��j^��>	�D<H�ԅ� �6�?�h��3��5ۭY��M�g��Kpc�Yg>��l��R�4���ƶf%��ج�U����M�`�
pIf� y��}ސ���/��6h�x*.��d�|���C�r �P�4�|�SEYW�������s�s=U`[W̾��`[��ܵp��I�8�pڛ����-��ÅN�n�i$ٚ%�H �|���N"�r�k��j��Dܚ��;�qdK�)�N�$�L�Yȇ�W�eG��ƕ���h��������^'hN�p��Q+�*@���m�5sp5k#q���c���puN��1��ޖ���7�Y�b�h#UJ�<���2>�X��������(�**���}o���|U��y~���C�*���ז��@w�5Y�$Q;�[���w�����-�R�P�C�v�|���4im����;�|��O��i�eK�Xq������"U�'�!�4�:�"_kl���\�R]�fo�.
`^�1otWB���FJቭ��N�q��[qv��H�17�M��A��E֎
�.�`����@��__��,4�}*2���N����M�|�ݰ$F:�������1�g�	���f�% ����&!)�h�s���7�
>G������#�!�!�ONy𚞙���H�卿p�����c�dW�<=[� Y^�ġ��`�;�4�1gx�YV� �y��x��S2�:TN^z��s��_(�=���|bgҗ��W���Ӵư͘~��U`)�y�h�Ǟc%�tPb�x�1��v-�Ig������봶w���d��d=$+�^��#^�kO���P'�̩�"Z%���4����vC'q�����,@����jp�1̇�MS8g��ւH]a�����V�&��`��a����>�����HW&��F>���as��p�F@%��l�,*��=g�}7�R�/7�k�!	��+��2y4�������T�y��,�y��~�����_���_A�aw��
�2T/��p�>AIV��ҡ��i��-Z�[LW�뎴��4�Zt~Z}[v�ĥm ?���^���l�`)�e9��t�1֬Q٧=UϾR+RG7��^�*�-�uL�<���{=�WX�0t{pDk��Q9�+bW]�-��_�T�&�d����pK��|S�@��U��4C��3f��N�sjL��Q���w�Q�)l�q����*r�c���)�t'�`��(�^��"�����8��r�k'4� P&�y�ك�c�J�8F/ч/��-2�`���O�e��c��Y&�I��g��fy��1!ڗ�/�Be��'g$5���BD��X^z�>&
�2,둱-�1GA�!��!�X�j,�G�$�oмΕ	\��v�S:�
f�Q���3D�}�|�&����K�I�9�>�Ner�!���y��Q���7�'�Z�\�~��koՐR}����Jv�a~��"A �Z��Vc(+�4Q���O�V,��x�л-��i�$la�j�W�azc03ęN��J��9����&E�ͧS��7�K�[����
K�ұ�VAU�J�J�u�C�v����d-���0
�k�� �tr�k+)�5�*�F}w[;�_R8TJn�� �����3�:->�A��������-
��%�a�q�ba:�,!ѧ�o���UQ�7@�����U����_zIx���BI �N�"�*^�}��pٿ��� ��i+�~S��%�T}�;�x��Us��ۀ�)Axs��:l�2�><B#"�>�q!m�{:DU�+�9x��R�ep ��� Q�Y���lv���8���pJ�GlA]�Rz#��j�&��6"K�p�m��^B+��:G�n�-��e��v��ߜ[G�)�m1f��t'�~12���{��Wt]%��e�n����o�W�D�
�J�u��Ӊ